
module top;

	reg p;

	inst #(15.99) ii0(p);

endmodule
