--* This source file is part of 'WAVES based' testbench.
--*   Copyright (C) ALDEC Inc.
--*
--* The IEEE Standard for Waveform and Vector Exchange to Support Design 
--*  and Test Verification (WAVES) is an formal notation inteneded for use 
--*  in all phases of the development of electronics system.  
--*
--* This VHDL file contains the declaration of the WAVES_GENERATOR package.
--
--  Title   : WAVES_GENERATOR
--
--  Library : This package shall be compiled into a current project library. 
--
--  Purpose : This package contains declaration of concurent procedure named WAVEFORM 
--            which generate - based on external Test Vector file - 
--            waveforms used as stimulus and outputs paterns 
--            for tested Unit Under Test (UUT).
--            This procedure is used in 'WAVES based' Test Bench 
--            automatically generated by Active VHDL Wizard.
--
-- --------------------------------------------------------------------
-- Modification history :
-- --------------------------------------------------------------------
--   Version:  1.0
--   Date   :  01 December 1997
--   Reason :  First version of 'WAVES based' Test Bench Wizard
-- --------------------------------------------------------------------

library IEEE;
use STD.textio.all;
use IEEE.waves_1164_frames.all;
use IEEE.waves_interface.all;
use work.waves_objects.all;
use work.uut_test_Pins.all;
use work.DESIGN_DECLARATIONS.all;

package WAVES_GENERATOR is
	procedure  WAVEFORM (
		signal WPL:			out WAVES_PORT_LIST; 
		signal END_VECTORS: 	out WAVES_TAG);
end WAVES_GENERATOR;

--------------------------------------------------------

package body WAVES_GENERATOR is

procedure WAVEFORM (
	signal WPL:			out WAVES_PORT_LIST; 
	signal END_VECTORS:	out WAVES_TAG) 
is

	variable vector: FILE_SLICE:= NEW_FILE_SLICE;
	
	type PINS_STIMULUS is array (TEST_PINS) of INTEGER;	
 
	procedure GET_MASK (
		ILINE: inout LINE; 
		variable POSITION_SET: inout PINS_STIMULUS) is
		
		variable POSITION: INTEGER;		
		variable DELTA: CHARACTER;
		variable GOOD: BOOLEAN:=TRUE;
	begin
		read (ILINE, DELTA); --skip @
		for PIN in POSITION_SET'range loop 
			read (ILINE, POSITION_SET(PIN));     
	   end loop;
	end;
		
	function SET_FRAME_TEMPLATE (STIMULATOR: INTEGER; STEP_TIME: DELAY_TIME; PIN: TEST_PINS) return FRAME_SET is
      variable WND: FRAME_SET;
      variable WINDOW_BEGIN, WINDOW_END: EVENT_TIME;
	begin
		if STIMULATOR = 1 then
			WND := NON_RETURN(STIM_BEGIN_DEFAULT);
		else
			WINDOW_BEGIN := WINDOW_TIME_LIST (PIN,START_T);
			WINDOW_END := WINDOW_TIME_LIST (PIN,END_T);
			if WINDOW_END = 0 ns then
				if STEP_TIME > 1 ps then
					WINDOW_END := STEP_TIME - 1 ps;
				else
					WINDOW_END := STEP_TIME;
				end if;					
			end if;
			
			WND := WINDOW(WINDOW_BEGIN, WINDOW_END);			
		end if;
		return WND;
	end;
      
	variable STIMULUS_SET: PINS_STIMULUS := (others=>1);
	variable PIN_TEMPLATE: FRAME_SET;
	variable PIN_FRAME: FRAME_DATA;
	variable PIN_MASK: PINSET:=NO_PINS;
	
	begin --of WAVEFORM procedure
		loop
			READ_FILE_SLICE (vector_file, VECTOR);  -- get first vector
			exit when vector.end_of_file;
			
			if VECTOR.TAG /= null then
				GET_MASK (VECTOR.TAG, STIMULUS_SET);       		
			end if;
			
			for PIN in STIMULUS_SET'range loop
				PIN_TEMPLATE := SET_FRAME_TEMPLATE(STIMULUS_SET(PIN), vector.fs_time, PIN);
				PIN_FRAME := BUILD_FRAME_DATA (( 1 => (+PIN, PIN_TEMPLATE)));
				PIN_MASK := NO_PINS;
				PIN_MASK(PIN) := TRUE;
				apply(WPL, VECTOR.codes.all, PIN_FRAME, PIN_MASK);
			end loop;
			
			delay (vector.fs_time);
		end loop;
		
		if VECTOR.TAG /= null then
			TAG (END_VECTORS, VECTOR.TAG.all);
		end if;
		
end WAVEFORM;
end WAVES_GENERATOR;
