--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:              4:59 PM, 4/20/99 *
--* Tested entity name:                             A8051_exp *
--* File name contains tested entity: $DSN\compile\A8051_exp.vhd *
--*************************************************************

library ieee;
use work.Types.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

	-- Add your library and packages declaration here ...

entity a8051_exp_tb is
end a8051_exp_tb;

architecture TB_ARCHITECTURE of a8051_exp_tb is
	-- Component declaration of the tested unit
	component A8051_exp
	port(
		CLK : in std_logic;
		KEY_0 : in std_logic;
		KEY_1 : in std_logic;
		KEY_2 : in std_logic;
		KEY_3 : in std_logic;
		KEY_4 : in std_logic;
		KEY_5 : in std_logic;
		KEY_6 : in std_logic;
		KEY_7 : in std_logic;
		KEY_8 : in std_logic;
		KEY_9 : in std_logic;
		RESET : in std_logic;
		nWRS : in std_logic;
		DATAS : in std_logic_vector(7 downto 0);
		BUSY : out std_logic;
		SCREEN : out ScrType );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal CLK : std_logic;
	signal KEY_0 : std_logic;
	signal KEY_1 : std_logic;
	signal KEY_2 : std_logic;
	signal KEY_3 : std_logic;
	signal KEY_4 : std_logic;
	signal KEY_5 : std_logic;
	signal KEY_6 : std_logic;
	signal KEY_7 : std_logic;
	signal KEY_8 : std_logic;
	signal KEY_9 : std_logic;
	signal RESET : std_logic;
	signal nWRS : std_logic;
	signal DATAS : std_logic_vector(7 downto 0):="00000000";
	-- Observed signals - signals mapped to the output ports of tested entity
	signal BUSY : std_logic;
	signal SCREEN : ScrType;

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : A8051_exp
		port map
			(CLK => CLK,
			KEY_0 => KEY_0,
			KEY_1 => KEY_1,
			KEY_2 => KEY_2,
			KEY_3 => KEY_3,
			KEY_4 => KEY_4,
			KEY_5 => KEY_5,
			KEY_6 => KEY_6,
			KEY_7 => KEY_7,
			KEY_8 => KEY_8,
			KEY_9 => KEY_9,
			RESET => RESET,
			nWRS => nWRS,
			DATAS => DATAS,
			BUSY => BUSY,
			SCREEN => SCREEN );

	--Below VHDL code is an inserted .\compile\keys.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

	KEY_0 <= '0';
	KEY_6 <= '0';
	nWRS <= '1';
	KEY_9 <= '0';
	KEY_8 <= '0';
	KEY_7 <= '0';
	KEY_5 <= '0';
	KEY_4 <= '0';
	KEY_3 <= '0';
	KEY_2 <= '0';
	KEY_1 <= '0';
    wait for 258100 ns; --0 ps
	nWRS <= '0';
    wait for 100 ns; --258100 ns
	nWRS <= '1';
    wait for 10900 ns; --258200 ns
	KEY_0 <= '1';
    wait for 200 ns; --269100 ns
	KEY_0 <= '0';
    wait for 99800 ns; --269300 ns
	nWRS <= '0';
    wait for 100 ns; --369100 ns
	nWRS <= '1';
    wait for 7800 ns; --369200 ns
	KEY_6 <= '1';
    wait for 500 ns; --377 us
	KEY_6 <= '0';
    wait for 222500 ns; --377500 ns
--	end of stimulus events
	wait;
end process; -- end of stimulus process
	
-- Add your stimulus here ...

DATA_CNT:
	process
	begin
		DATAS<=DATAS + "00000001";
		wait for 300 ns;	
	end process;
	
RST_CRC: process
          begin
          	RESET<='1';
          	wait for 1 us;
          	RESET<='0';
          	wait;
          end process;           

 CLK_GEN: process
		  begin
				CLK<= '1';
		  		wait for 0.01 us;
		  		CLK<= '0';
		  		wait for 0.01 us;
		  end process;	

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_A8051_exp of a8051_exp_tb is
	for TB_ARCHITECTURE
		for UUT : A8051_exp
			use entity work.A8051_exp(A8051_exp);
		end for;
	end for;
end TESTBENCH_FOR_A8051_exp;

