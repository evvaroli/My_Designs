library ieee;
use ieee.std_logic_1164.all;

package twos_complement_types is

  type twos_complement is array (natural range <>) of std_ulogic;

end twos_complement_types;
