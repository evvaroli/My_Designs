
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity player_font is
	port (
		angle: in STD_LOGIC_VECTOR (1 downto 0);
		addr: in STD_LOGIC_VECTOR (5 downto 0);
		M: out STD_LOGIC_VECTOR (0 to 31)
		);
end player_font;

architecture player_font of player_font is
	type rom_array is array (NATURAL range <>)  
	of STD_LOGIC_VECTOR (0 to 31);
	constant rom1: rom_array := (
	"11110000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"11000000000000000000000000000000",
	"11000000000000000000000000000000"
	);
begin
	process(addr)
	variable j: integer;				
	begin 
		j := conv_integer(addr);
			M <= rom1(j);
	end process; 
end player_font;