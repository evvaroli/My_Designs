// (c) Aldec, Inc.
// All rights reserved.
//
// Last modified: $Date: 2009-09-03 16:57:08 +0200 (Thu, 03 Sep 2009) $
// $Revision: 121928 $


// ROM : 256 8-bit words - multiplication with c3=8 coefficient
module rom_rtl_c3(
				input [7:0] addr,
				output reg [15:0] data
				);


always @(addr)
begin
	case (addr)
		8'd0   : data = 11'd0;
		8'd1   : data = 11'd8;
		8'd2   : data = 11'd16;
		8'd3   : data = 11'd24;
		8'd4   : data = 11'd32;
		8'd5   : data = 11'd40;
		8'd6   : data = 11'd48;
		8'd7   : data = 11'd56;
		8'd8   : data = 11'd64;
		8'd9   : data = 11'd72;
		8'd10  : data = 11'd80;
		8'd11  : data = 11'd88;
		8'd12  : data = 11'd96;
		8'd13  : data = 11'd104;
		8'd14  : data = 11'd112;
		8'd15  : data = 11'd120;
		8'd16  : data = 11'd128;
		8'd17  : data = 11'd136;
		8'd18  : data = 11'd144;
		8'd19  : data = 11'd152;
		8'd20  : data = 11'd160;
		8'd21  : data = 11'd168;
		8'd22  : data = 11'd176;
		8'd23  : data = 11'd184;
		8'd24  : data = 11'd192;
		8'd25  : data = 11'd200;
		8'd26  : data = 11'd208;
		8'd27  : data = 11'd216;
		8'd28  : data = 11'd224;
		8'd29  : data = 11'd232;
		8'd30  : data = 11'd240;
		8'd31  : data = 11'd248;
		8'd32  : data = 11'd256;
		8'd33  : data = 11'd264;
		8'd34  : data = 11'd272;
		8'd35  : data = 11'd280;
		8'd36  : data = 11'd288;
		8'd37  : data = 11'd296;
		8'd38  : data = 11'd304;
		8'd39  : data = 11'd312;
		8'd40  : data = 11'd320;
		8'd41  : data = 11'd328;
		8'd42  : data = 11'd336;
		8'd43  : data = 11'd344;
		8'd44  : data = 11'd352;
		8'd45  : data = 11'd360;
		8'd46  : data = 11'd368;
		8'd47  : data = 11'd376;
		8'd48  : data = 11'd384;
		8'd49  : data = 11'd392;
		8'd50  : data = 11'd400;
		8'd51  : data = 11'd408;
		8'd52  : data = 11'd416;
		8'd53  : data = 11'd424;
		8'd54  : data = 11'd432;
		8'd55  : data = 11'd440;
		8'd56  : data = 11'd448;
		8'd57  : data = 11'd456;
		8'd58  : data = 11'd464;
		8'd59  : data = 11'd472;
		8'd60  : data = 11'd480;
		8'd61  : data = 11'd488;
		8'd62  : data = 11'd496;
		8'd63  : data = 11'd504;
		8'd64  : data = 11'd512;
		8'd65  : data = 11'd520;
		8'd66  : data = 11'd528;
		8'd67  : data = 11'd536;
		8'd68  : data = 11'd544;
		8'd69  : data = 11'd552;
		8'd70  : data = 11'd560;
		8'd71  : data = 11'd568;
		8'd72  : data = 11'd576;
		8'd73  : data = 11'd584;
		8'd74  : data = 11'd592;
		8'd75  : data = 11'd600;
		8'd76  : data = 11'd608;
		8'd77  : data = 11'd616;
		8'd78  : data = 11'd624;
		8'd79  : data = 11'd632;
		8'd80  : data = 11'd640;
		8'd81  : data = 11'd648;
		8'd82  : data = 11'd656;
		8'd83  : data = 11'd664;
		8'd84  : data = 11'd672;
		8'd85  : data = 11'd680;
		8'd86  : data = 11'd688;
		8'd87  : data = 11'd696;
		8'd88  : data = 11'd704;
		8'd89  : data = 11'd712;
		8'd90  : data = 11'd720;
		8'd91  : data = 11'd728;
		8'd92  : data = 11'd736;
		8'd93  : data = 11'd744;
		8'd94  : data = 11'd752;
		8'd95  : data = 11'd760;
		8'd96  : data = 11'd768;
		8'd97  : data = 11'd776;
		8'd98  : data = 11'd784;
		8'd99  : data = 11'd792;
		8'd100 : data = 11'd800;
		8'd101 : data = 11'd808;
		8'd102 : data = 11'd816;
		8'd103 : data = 11'd824;
		8'd104 : data = 11'd832;
		8'd105 : data = 11'd840;
		8'd106 : data = 11'd848;
		8'd107 : data = 11'd856;
		8'd108 : data = 11'd864;
		8'd109 : data = 11'd872;
		8'd110 : data = 11'd880;
		8'd111 : data = 11'd888;
		8'd112 : data = 11'd896;
		8'd113 : data = 11'd904;
		8'd114 : data = 11'd912;
		8'd115 : data = 11'd920;
		8'd116 : data = 11'd928;
		8'd117 : data = 11'd936;
		8'd118 : data = 11'd944;
		8'd119 : data = 11'd952;
		8'd120 : data = 11'd960;
		8'd121 : data = 11'd968;
		8'd122 : data = 11'd976;
		8'd123 : data = 11'd984;
		8'd124 : data = 11'd992;
		8'd125 : data = 11'd1000;
		8'd126 : data = 11'd1008;
		8'd127 : data = 11'd1016;
		8'd128 : data = 11'd1024;
		8'd129 : data = 11'd1032;
		8'd130 : data = 11'd1040;
		8'd131 : data = 11'd1048;
		8'd132 : data = 11'd1056;
		8'd133 : data = 11'd1064;
		8'd134 : data = 11'd1072;
		8'd135 : data = 11'd1080;
		8'd136 : data = 11'd1088;
		8'd137 : data = 11'd1096;
		8'd138 : data = 11'd1104;
		8'd139 : data = 11'd1112;
		8'd140 : data = 11'd1120;
		8'd141 : data = 11'd1128;
		8'd142 : data = 11'd1136;
		8'd143 : data = 11'd1144;
		8'd144 : data = 11'd1152;
		8'd145 : data = 11'd1160;
		8'd146 : data = 11'd1168;
		8'd147 : data = 11'd1176;
		8'd148 : data = 11'd1184;
		8'd149 : data = 11'd1192;
		8'd150 : data = 11'd1200;
		8'd151 : data = 11'd1208;
		8'd152 : data = 11'd1216;
		8'd153 : data = 11'd1224;
		8'd154 : data = 11'd1232;
		8'd155 : data = 11'd1240;
		8'd156 : data = 11'd1248;
		8'd157 : data = 11'd1256;
		8'd158 : data = 11'd1264;
		8'd159 : data = 11'd1272;
		8'd160 : data = 11'd1280;
		8'd161 : data = 11'd1288;
		8'd162 : data = 11'd1296;
		8'd163 : data = 11'd1304;
		8'd164 : data = 11'd1312;
		8'd165 : data = 11'd1320;
		8'd166 : data = 11'd1328;
		8'd167 : data = 11'd1336;
		8'd168 : data = 11'd1344;
		8'd169 : data = 11'd1352;
		8'd170 : data = 11'd1360;
		8'd171 : data = 11'd1368;
		8'd172 : data = 11'd1376;
		8'd173 : data = 11'd1384;
		8'd174 : data = 11'd1392;
		8'd175 : data = 11'd1400;
		8'd176 : data = 11'd1408;
		8'd177 : data = 11'd1416;
		8'd178 : data = 11'd1424;
		8'd179 : data = 11'd1432;
		8'd180 : data = 11'd1440;
		8'd181 : data = 11'd1448;
		8'd182 : data = 11'd1456;
		8'd183 : data = 11'd1464;
		8'd184 : data = 11'd1472;
		8'd185 : data = 11'd1480;
		8'd186 : data = 11'd1488;
		8'd187 : data = 11'd1496;
		8'd188 : data = 11'd1504;
		8'd189 : data = 11'd1512;
		8'd190 : data = 11'd1520;
		8'd191 : data = 11'd1528;
		8'd192 : data = 11'd1536;
		8'd193 : data = 11'd1544;
		8'd194 : data = 11'd1552;
		8'd195 : data = 11'd1560;
		8'd196 : data = 11'd1568;
		8'd197 : data = 11'd1576;
		8'd198 : data = 11'd1584;
		8'd199 : data = 11'd1592;
		8'd200 : data = 11'd1600;
		8'd201 : data = 11'd1608;
		8'd202 : data = 11'd1616;
		8'd203 : data = 11'd1624;
		8'd204 : data = 11'd1632;
		8'd205 : data = 11'd1640;
		8'd206 : data = 11'd1648;
		8'd207 : data = 11'd1656;
		8'd208 : data = 11'd1664;
		8'd209 : data = 11'd1672;
		8'd210 : data = 11'd1680;
		8'd211 : data = 11'd1688;
		8'd212 : data = 11'd1696;
		8'd213 : data = 11'd1704;
		8'd214 : data = 11'd1712;
		8'd215 : data = 11'd1720;
		8'd216 : data = 11'd1728;
		8'd217 : data = 11'd1736;
		8'd218 : data = 11'd1744;
		8'd219 : data = 11'd1752;
		8'd220 : data = 11'd1760;
		8'd221 : data = 11'd1768;
		8'd222 : data = 11'd1776;
		8'd223 : data = 11'd1784;
		8'd224 : data = 11'd1792;
		8'd225 : data = 11'd1800;
		8'd226 : data = 11'd1808;
		8'd227 : data = 11'd1816;
		8'd228 : data = 11'd1824;
		8'd229 : data = 11'd1832;
		8'd230 : data = 11'd1840;
		8'd231 : data = 11'd1848;
		8'd232 : data = 11'd1856;
		8'd233 : data = 11'd1864;
		8'd234 : data = 11'd1872;
		8'd235 : data = 11'd1880;
		8'd236 : data = 11'd1888;
		8'd237 : data = 11'd1896;
		8'd238 : data = 11'd1904;
		8'd239 : data = 11'd1912;
		8'd240 : data = 11'd1920;
		8'd241 : data = 11'd1928;
		8'd242 : data = 11'd1936;
		8'd243 : data = 11'd1944;
		8'd244 : data = 11'd1952;
		8'd245 : data = 11'd1960;
		8'd246 : data = 11'd1968;
		8'd247 : data = 11'd1976;
		8'd248 : data = 11'd1984;
		8'd249 : data = 11'd1992;
		8'd250 : data = 11'd2000;
		8'd251 : data = 11'd2008;
		8'd252 : data = 11'd2016;
		8'd253 : data = 11'd2024;
		8'd254 : data = 11'd2032;
		8'd255 : data = 11'd2040;
    endcase
end

endmodule
