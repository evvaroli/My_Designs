`timescale 1ns/1ps
module tb;

logic clk,rst;
logic [7:0] in,out;

initial begin 
	rst = 1;
	clk = 0;
	#10;
	rst = 0;
end

always #5 clk = ~clk;

fir dut(
	.clk(clk),
	.rst(rst),
	.inp(in),
	.outp(out));

initial begin
	in = 8'b10010010;
    #10; //0
	in = 8'b01000000;
    #10; //10000
	in = 8'b00000100;
    #10; //20000
	in = 8'b00110001;
    #10; //30000
	in = 8'b10000110;
    #10; //40000
	in = 8'b11000110;
    #10; //50000
	in = 8'b00110010;
    #10; //60000
	in = 8'b00001001;
    #10; //70000
	in = 8'b10000000;
    #10; //80000
	in = 8'b10000110;
    #10; //90000
	in = 8'b10111011;
    #10; //100000
	in = 8'b10011110;
    #10; //110000
	in = 8'b11110110;
    #10; //120000
	in = 8'b11000110;
    #10; //130000
	in = 8'b11111100;
    #10; //140000
	in = 8'b01100011;
    #10; //150000
	in = 8'b01100010;
    #10; //160000
	in = 8'b01010101;
    #10; //170000
	in = 8'b11110010;
    #10; //180000
	in = 8'b00111011;
    #10; //190000
	in = 8'b00001001;
    #10; //200000
	in = 8'b11000111;
    #10; //210000
	in = 8'b11111001;
    #10; //220000
	in = 8'b01100111;
    #10; //230000
	in = 8'b01110100;
    #10; //240000
	in = 8'b01100010;
    #10; //250000
	in = 8'b10101110;
    #10; //260000
	in = 8'b01011110;
    #10; //270000
	in = 8'b00010110;
    #10; //280000
	in = 8'b00110010;
    #10; //290000
	in = 8'b00110001;
	#10;
	$finish;
end

endmodule : tb
