library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity title_prom is
    port (
        addr: in STD_LOGIC_VECTOR (3 downto 0);
        M: out STD_LOGIC_VECTOR (0 to 31)
    );
end title_prom;

architecture title_prom of title_prom is
type rom_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 31);	
constant rom: rom_array := (
	"01111110000011000001101000000010", 		--0
	"01000001000011000001101000000010", 		--1
	"01000000100010100010101000000010", 		--2
	"01000000010010100010101000000010", 		--3
	"01000000001010100010101000000010", 		--4
	"01000000001010010100101000000010", 		--5
	"01000000001010010100101000000010", 		--6
	"01000000001010010100101111111110", 		--7
	"01000000001010001000101000000010", 		--8
	"01000000001010001000101000000010", 		--9
	"01000000001010001000101000000010", 		--10
	"01000000001010000000101000000010", 		--11
	"01000000010010000000101000000010", 		--12
	"01000000100010000000101000000010", 		--13
	"01000001000010000000101000000010", 		--14
	"01111110000010000000101000000010"	 		--15
	);				   
	
	begin
	
	  process(addr)
	  variable j: integer;
	  begin 
	    j := conv_integer(addr);
	    M <= rom(j);
	  end process;
 
end title_prom;