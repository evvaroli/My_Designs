
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity tank_sprite is
	port (
		angle: in STD_LOGIC_VECTOR(1 downto 0);
		addr: in STD_LOGIC_VECTOR (5 downto 0);
		M: out STD_LOGIC_VECTOR (0 to 31)
		);
end tank_sprite;

architecture tank_sprite of tank_sprite is
	type rom_array is array (NATURAL range <>)  
	of STD_LOGIC_VECTOR (0 to 31);
	
	constant rom1: rom_array:= (
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000011111110000000000000",
	"00000000001100000001000000000000",
	"00000000010000000000100000000000",
	"00000000100000000000100000000000",
	"00011111100000000000111111111111",
	"01100000100000000000100000001001",
	"10001111100011111111100000001001",
	"10010000101100000000100000001001",
	"11110000110000000000010000001111",
	"11110000100000000000011111111100",
	"11111111100000000000001111111100",
	"11110000100000000000001100001100",
	"11111111111000000000111100001100",
	"11111111111100111111111100001100",
	"11100000011111000001111111111000",
	"10000000010001101111000000001000",
	"10011011110001010001000000000100",
	"11100100001111111111111011110100",
	"10000100000000000000000100001100",
	"10000100000000000000000100000100",
	"10000100000000000000000100000100",
	"11111111111111111111111111111100",
	"10111111111111111111111111111100",
	"01111111111111111111111111101000",
	"01010010010010010010010011011000",
	"00101001001001001001001001110000",
	"00111111111111111111111111000000"
	);	  
	
	constant rom2: rom_array := (
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000011111110000000001100",
	"00000000001100000001000000110010",
	"00000000010000000000100011010010",
	"00000000100000000000101100011001",
	"00011111100000000000110000001001",
	"01100000100000000000100000001110",
	"10001111100011111111100000011000",
	"10010000101100000000100001111000",
	"11110000110000000000010110001000",
	"11110000100000000000011111111100",
	"11111111100000000000001111111100",
	"11110000100000000000001100001100",
	"11111111111000000000111100001100",
	"11111111111100111111111100001100",
	"11100000011111000001111111111000",
	"10000000010001101111000000001000",
	"10011011110001010001000000000100",
	"11100100001111111111111011110100",
	"10000100000000000000000100001100",
	"10000100000000000000000100000100",
	"10000100000000000000000100000100",
	"11111111111111111111111111111100",
	"10111111111111111111111111111100",
	"01111111111111111111111111101000",
	"01010010010010010010010011011000",
	"00101001001001001001001001110000",
	"00111111111111111111111111000000"
	);
	constant rom3: rom_array := (
	"00000000000000000000000000010000",
	"00000000000000000000000000101000",
	"00000000000011111110000011000100",
	"00000000001100000001000101100010",
	"00000000010000000000101000110100",
	"00000000100000000000110000011000",
	"00011111100000000000100000001000",
	"01100000100000000000100000010000",
	"10001111100011111111100000110000",
	"10010000101100000000100001111000",
	"11110000110000000000010010001100",
	"11110000100000000000010111111100",
	"11111111100000000000001111111100",
	"11110000100000000000001100001100",
	"11111111111000000000111100001100",
	"11111111111100111111111100001100",
	"11100000011111000001111111111000",
	"10000000010001101111000000001000",
	"10011011110001010001000000000100",
	"11100100001111111111111011110100",
	"10000100000000000000000100001100",
	"10000100000000000000000100000100",
	"10000100000000000000000100000100",
	"11111111111111111111111111111100",
	"10111111111111111111111111111100",
	"01111111111111111111111111101000",
	"01010010010010010010010011011000",
	"00101001001001001001001001110000",
	"00111111111111111111111111000000"
	);
begin
	process(addr)
		variable j: integer;	
	begin
		j := conv_integer(addr);
		if angle = "00" then
			M <= rom1(j);
		elsif angle = "11" then
			M <= rom3(j);
		else
			M <= rom2(j);
		end if;
	end process; 
end tank_sprite;