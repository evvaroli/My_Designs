
module top;

	reg p;

	inst #(15) ii0(p);

endmodule
