module AND2 (A0, A1, Y);

input A0;
wire A0;
input A1;
wire A1;
output Y;
wire Y;

// add your declarations here

// add your code here
	assign Y = A0 & A1;
endmodule 
