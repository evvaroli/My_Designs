-- Copyright (c) Aldec, Inc.
-- All rights reserved.
--
-- Last modified: $Date: 2007-11-29 17:49:29 +0100 (Thu, 29 Nov 2007) $
-- $Revision: 70682 $

entity tb is
end entity;
