
`timescale 1ps / 1ps
module filter_tb;


//Internal signals declarations:
reg [3:0]NI;
reg CLK;
reg RESET;
wire [3:0]NO;

//---
integer res_file;
								  
initial
begin
	res_file = $fopen ("results_verlog.txt");
end	

always @ (NI or NO or CLK or RESET)
begin
	$fdisplay (res_file, " %d ps %b %b %b %b", $time,
				NI, NO, CLK, RESET);
end

//--

// Unit Under Test port map
	filter UUT (
		.NI(NI),
		.CLK(CLK),
		.RESET(RESET),
		.NO(NO));

initial
	$monitor($realtime,,"ps %h %h %h %h ",NI,CLK,RESET,NO);


initial
begin : STIMUL // begin of stimulus process
	#0
	NI = 4'b0001;
	CLK = 1'b0;
	RESET = 1'b1;
    #10000; //0
	CLK = 1'b1;
    #10000; //10000
	CLK = 1'b0;
    #10000; //20000
	CLK = 1'b1;
    #10000; //30000
	CLK = 1'b0;
    #5000; //40000
	RESET = 1'b0;
    #5000; //45000
	CLK = 1'b1;
    #10000; //50000
	CLK = 1'b0;
    #10000; //60000
	CLK = 1'b1;
    #10000; //70000
	CLK = 1'b0;
    #10000; //80000
	CLK = 1'b1;
    #10000; //90000
	CLK = 1'b0;
    #10000; //100000
	CLK = 1'b1;
    #10000; //110000
	CLK = 1'b0;
    #10000; //120000
	CLK = 1'b1;
    #10000; //130000
	CLK = 1'b0;
    #10000; //140000
	CLK = 1'b1;
    #10000; //150000
	CLK = 1'b0;
    #10000; //160000
	CLK = 1'b1;
    #10000; //170000
	CLK = 1'b0;
    #10000; //180000
	CLK = 1'b1;
    #10000; //190000
	CLK = 1'b0;
    #10000; //200000
	CLK = 1'b1;
    #10000; //210000
	CLK = 1'b0;
    #10000; //220000
	CLK = 1'b1;
    #10000; //230000
	CLK = 1'b0;
    #10000; //240000
	CLK = 1'b1;
    #10000; //250000
	CLK = 1'b0;
    #10000; //260000
	CLK = 1'b1;
    #10000; //270000
	CLK = 1'b0;
    #10000; //280000
	CLK = 1'b1;
    #10000; //290000
	CLK = 1'b0;
    #10000; //300000
	CLK = 1'b1;
    #10000; //310000
	CLK = 1'b0;
    #10000; //320000
	CLK = 1'b1;
    #10000; //330000
	CLK = 1'b0;
    #10000; //340000
	CLK = 1'b1;
    #10000; //350000
	CLK = 1'b0;
    #10000; //360000
	CLK = 1'b1;
    #10000; //370000
	CLK = 1'b0;
    #10000; //380000
	CLK = 1'b1;
    #10000; //390000
	CLK = 1'b0;
    #10000; //400000
	CLK = 1'b1;
    #10000; //410000
	CLK = 1'b0;
    #10000; //420000
	CLK = 1'b1;
    #10000; //430000
	CLK = 1'b0;
    #10000; //440000
	CLK = 1'b1;
    #10000; //450000
	CLK = 1'b0;
    #10000; //460000
	CLK = 1'b1;
    #10000; //470000
	CLK = 1'b0;
    #10000; //480000
	CLK = 1'b1;
    #10000; //490000
	CLK = 1'b0;
    #10000; //500000
	CLK = 1'b1;
    #10000; //510000
	CLK = 1'b0;
    #10000; //520000
	CLK = 1'b1;
    #10000; //530000
	CLK = 1'b0;
    #10000; //540000
	CLK = 1'b1;
    #10000; //550000
	CLK = 1'b0;
    #10000; //560000
	CLK = 1'b1;
    #10000; //570000
	CLK = 1'b0;
    #10000; //580000
	CLK = 1'b1;
    #10000; //590000
	CLK = 1'b0;
    #10000; //600000
	CLK = 1'b1;
    #10000; //610000
	CLK = 1'b0;
    #10000; //620000
	CLK = 1'b1;
    #10000; //630000
	CLK = 1'b0;
    #10000; //640000
	CLK = 1'b1;
    #10000; //650000
	CLK = 1'b0;
    #10000; //660000
	CLK = 1'b1;
    #10000; //670000
	CLK = 1'b0;
    #10000; //680000
	CLK = 1'b1;
    #10000; //690000
	CLK = 1'b0;
    #10000; //700000
	CLK = 1'b1;
    #10000; //710000
	CLK = 1'b0;
    #10000; //720000
	CLK = 1'b1;
    #10000; //730000
	CLK = 1'b0;
    #10000; //740000
	CLK = 1'b1;
    #10000; //750000
	CLK = 1'b0;
    #10000; //760000
	CLK = 1'b1;
    #10000; //770000
	CLK = 1'b0;
    #10000; //780000
	CLK = 1'b1;
    #10000; //790000
	CLK = 1'b0;
    #10000; //800000
	CLK = 1'b1;
    #10000; //810000
	CLK = 1'b0;
    #10000; //820000
	CLK = 1'b1;
    #10000; //830000
	CLK = 1'b0;
    #10000; //840000
	CLK = 1'b1;
    #10000; //850000
	CLK = 1'b0;
    #10000; //860000
	CLK = 1'b1;
    #10000; //870000
	CLK = 1'b0;
    #10000; //880000
	CLK = 1'b1;
    #10000; //890000
	CLK = 1'b0;
    #10000; //900000
	CLK = 1'b1;
    #10000; //910000
	CLK = 1'b0;
    #10000; //920000
	CLK = 1'b1;
    #10000; //930000
	CLK = 1'b0;
    #10000; //940000
	CLK = 1'b1;
    #10000; //950000
	CLK = 1'b0;
    #10000; //960000
	CLK = 1'b1;
    #10000; //970000
	CLK = 1'b0;
    #10000; //980000
	CLK = 1'b1;
    #10000; //990000
	CLK = 1'b0;
    #10000; //1000000
	CLK = 1'b1;
    #10000; //1010000
	CLK = 1'b0;
    #10000; //1020000
	CLK = 1'b1;
    #10000; //1030000
	CLK = 1'b0;
    #10000; //1040000
	CLK = 1'b1;
    #10000; //1050000
	CLK = 1'b0;
    #10000; //1060000
	CLK = 1'b1;
    #10000; //1070000
	CLK = 1'b0;
    #10000; //1080000
	CLK = 1'b1;
    #10000; //1090000
	CLK = 1'b0;
    #10000; //1100000
	CLK = 1'b1;
    #10000; //1110000
	CLK = 1'b0;
    #10000; //1120000
	CLK = 1'b1;
    #10000; //1130000
	CLK = 1'b0;
    #10000; //1140000
	CLK = 1'b1;
    #10000; //1150000
	CLK = 1'b0;
    #10000; //1160000
	CLK = 1'b1;
    #10000; //1170000
	CLK = 1'b0;
    #10000; //1180000
	CLK = 1'b1;
    #10000; //1190000
	CLK = 1'b0;
    #10000; //1200000
	CLK = 1'b1;
    #10000; //1210000
	CLK = 1'b0;
    #10000; //1220000
	CLK = 1'b1;
    #10000; //1230000
	CLK = 1'b0;
    #10000; //1240000
	CLK = 1'b1;
    #10000; //1250000
	CLK = 1'b0;
    #10000; //1260000
	CLK = 1'b1;
    #10000; //1270000
	CLK = 1'b0;
    #10000; //1280000
	CLK = 1'b1;
    #10000; //1290000
	CLK = 1'b0;
    #10000; //1300000
	CLK = 1'b1;
    #10000; //1310000
	CLK = 1'b0;
    #10000; //1320000
	CLK = 1'b1;
    #10000; //1330000
	CLK = 1'b0;
    #10000; //1340000
	CLK = 1'b1;
    #10000; //1350000
	CLK = 1'b0;
    #10000; //1360000
	CLK = 1'b1;
    #10000; //1370000
	CLK = 1'b0;
    #10000; //1380000
	CLK = 1'b1;
    #10000; //1390000
	CLK = 1'b0;
    #10000; //1400000
	CLK = 1'b1;
    #10000; //1410000
	CLK = 1'b0;
    #10000; //1420000
	CLK = 1'b1;
    #10000; //1430000
	CLK = 1'b0;
    #10000; //1440000
	CLK = 1'b1;
    #10000; //1450000
	CLK = 1'b0;
    #10000; //1460000
	CLK = 1'b1;
    #10000; //1470000
	CLK = 1'b0;
    #10000; //1480000
	CLK = 1'b1;
    #10000; //1490000
	CLK = 1'b0;
    #10000; //1500000
	CLK = 1'b1;
    #10000; //1510000
	CLK = 1'b0;
    #10000; //1520000
	CLK = 1'b1;
    #10000; //1530000
	CLK = 1'b0;
    #10000; //1540000
	CLK = 1'b1;
    #10000; //1550000
	CLK = 1'b0;
    #10000; //1560000
	CLK = 1'b1;
    #10000; //1570000
	CLK = 1'b0;
    #10000; //1580000
	CLK = 1'b1;
    #10000; //1590000
	CLK = 1'b0;
    #10000; //1600000
	CLK = 1'b1;
    #10000; //1610000
	CLK = 1'b0;
    #10000; //1620000
	CLK = 1'b1;
    #10000; //1630000
	CLK = 1'b0;
    #10000; //1640000
	CLK = 1'b1;
    #10000; //1650000
	CLK = 1'b0;
    #10000; //1660000
	CLK = 1'b1;
    #10000; //1670000
	CLK = 1'b0;
    #10000; //1680000
	CLK = 1'b1;
    #10000; //1690000
	CLK = 1'b0;
    #10000; //1700000
	CLK = 1'b1;
    #10000; //1710000
	CLK = 1'b0;
    #10000; //1720000
	CLK = 1'b1;
    #10000; //1730000
	CLK = 1'b0;
    #10000; //1740000
	CLK = 1'b1;
    #10000; //1750000
	CLK = 1'b0;
    #10000; //1760000
	CLK = 1'b1;
    #10000; //1770000
	CLK = 1'b0;
    #10000; //1780000
	CLK = 1'b1;
    #10000; //1790000
	CLK = 1'b0;
    #10000; //1800000
	CLK = 1'b1;
    #10000; //1810000
	CLK = 1'b0;
    #10000; //1820000
	CLK = 1'b1;
    #10000; //1830000
	CLK = 1'b0;
    #10000; //1840000
	CLK = 1'b1;
    #10000; //1850000
	CLK = 1'b0;
    #10000; //1860000
	CLK = 1'b1;
    #10000; //1870000
	CLK = 1'b0;
    #10000; //1880000
	CLK = 1'b1;
    #10000; //1890000
	CLK = 1'b0;
    #10000; //1900000
	CLK = 1'b1;
    #10000; //1910000
	CLK = 1'b0;
    #10000; //1920000
	CLK = 1'b1;
    #10000; //1930000
	CLK = 1'b0;
    #10000; //1940000
	CLK = 1'b1;
    #10000; //1950000
	CLK = 1'b0;
    #10000; //1960000
	CLK = 1'b1;
    #10000; //1970000
	CLK = 1'b0;
    #10000; //1980000
	CLK = 1'b1;
    #10000; //1990000
	CLK = 1'b0;
    #10000; //2000000
	CLK = 1'b1;
    #10000; //2010000
	CLK = 1'b0;
    #10000; //2020000
	CLK = 1'b1;
    #10000; //2030000
	CLK = 1'b0;
    #10000; //2040000
	CLK = 1'b1;
    #10000; //2050000
	CLK = 1'b0;
    #10000; //2060000
	CLK = 1'b1;
    #10000; //2070000
	CLK = 1'b0;
    #10000; //2080000
	CLK = 1'b1;
    #10000; //2090000
	CLK = 1'b0;
    #10000; //2100000
	CLK = 1'b1;
    #10000; //2110000
	CLK = 1'b0;
    #10000; //2120000
	CLK = 1'b1;
    #10000; //2130000
	CLK = 1'b0;
    #5000; //2140000
	NI = 4'b1111;
    #5000; //2145000
	CLK = 1'b1;
    #10000; //2150000
	CLK = 1'b0;
    #10000; //2160000
	CLK = 1'b1;
    #10000; //2170000
	CLK = 1'b0;
    #10000; //2180000
	CLK = 1'b1;
    #10000; //2190000
	CLK = 1'b0;
    #10000; //2200000
	CLK = 1'b1;
    #10000; //2210000
	CLK = 1'b0;
    #10000; //2220000
	CLK = 1'b1;
    #10000; //2230000
	CLK = 1'b0;
    #10000; //2240000
	CLK = 1'b1;
    #10000; //2250000
	CLK = 1'b0;
    #10000; //2260000
	CLK = 1'b1;
    #10000; //2270000
	CLK = 1'b0;
    #10000; //2280000
	CLK = 1'b1;
    #10000; //2290000
	CLK = 1'b0;
    #10000; //2300000
	CLK = 1'b1;
    #10000; //2310000
	CLK = 1'b0;
    #10000; //2320000
	CLK = 1'b1;
    #10000; //2330000
	CLK = 1'b0;
    #10000; //2340000
	CLK = 1'b1;
    #10000; //2350000
	CLK = 1'b0;
    #10000; //2360000
	CLK = 1'b1;
    #10000; //2370000
	CLK = 1'b0;
    #10000; //2380000
	CLK = 1'b1;
    #10000; //2390000
	CLK = 1'b0;
    #10000; //2400000
	CLK = 1'b1;
    #10000; //2410000
	CLK = 1'b0;
    #10000; //2420000
	CLK = 1'b1;
    #10000; //2430000
	CLK = 1'b0;
    #10000; //2440000
	CLK = 1'b1;
    #10000; //2450000
	CLK = 1'b0;
    #10000; //2460000
	CLK = 1'b1;
    #10000; //2470000
	CLK = 1'b0;
    #10000; //2480000
	CLK = 1'b1;
    #10000; //2490000
	CLK = 1'b0;
    #10000; //2500000
	CLK = 1'b1;
    #10000; //2510000
	CLK = 1'b0;
    #10000; //2520000
	CLK = 1'b1;
    #10000; //2530000
	CLK = 1'b0;
    #10000; //2540000
	CLK = 1'b1;
    #10000; //2550000
	CLK = 1'b0;
    #10000; //2560000
	CLK = 1'b1;
    #10000; //2570000
	CLK = 1'b0;
    #10000; //2580000
	CLK = 1'b1;
    #10000; //2590000
	CLK = 1'b0;
    #10000; //2600000
	CLK = 1'b1;
    #10000; //2610000
	CLK = 1'b0;
    #10000; //2620000
	CLK = 1'b1;
    #10000; //2630000
	CLK = 1'b0;
    #10000; //2640000
	CLK = 1'b1;
    #10000; //2650000
	CLK = 1'b0;
    #10000; //2660000
	CLK = 1'b1;
    #10000; //2670000
	CLK = 1'b0;
    #10000; //2680000
	CLK = 1'b1;
    #10000; //2690000
	CLK = 1'b0;
    #10000; //2700000
	CLK = 1'b1;
    #10000; //2710000
	CLK = 1'b0;
    #10000; //2720000
	CLK = 1'b1;
    #10000; //2730000
	CLK = 1'b0;
    #10000; //2740000
	CLK = 1'b1;
    #10000; //2750000
	CLK = 1'b0;
    #10000; //2760000
	CLK = 1'b1;
    #10000; //2770000
	CLK = 1'b0;
    #10000; //2780000
	CLK = 1'b1;
    #10000; //2790000
	CLK = 1'b0;
    #10000; //2800000
	CLK = 1'b1;
    #10000; //2810000
	CLK = 1'b0;
    #10000; //2820000
	CLK = 1'b1;
    #10000; //2830000
	CLK = 1'b0;
    #10000; //2840000
	CLK = 1'b1;
    #10000; //2850000
	CLK = 1'b0;
    #10000; //2860000
	CLK = 1'b1;
    #10000; //2870000
	CLK = 1'b0;
    #10000; //2880000
	CLK = 1'b1;
    #10000; //2890000
	CLK = 1'b0;
    #10000; //2900000
	CLK = 1'b1;
    #10000; //2910000
	CLK = 1'b0;
    #10000; //2920000
	CLK = 1'b1;
    #10000; //2930000
	CLK = 1'b0;
    #10000; //2940000
	CLK = 1'b1;
    #10000; //2950000
	CLK = 1'b0;
    #10000; //2960000
	CLK = 1'b1;
    #10000; //2970000
	CLK = 1'b0;
    #10000; //2980000
	CLK = 1'b1;
    #10000; //2990000
	CLK = 1'b0;
    #10000; //3000000
	CLK = 1'b1;
    #10000; //3010000
	CLK = 1'b0;
    #10000; //3020000
	CLK = 1'b1;
    #10000; //3030000
	CLK = 1'b0;
    #10000; //3040000
	CLK = 1'b1;
    #10000; //3050000
	CLK = 1'b0;
    #10000; //3060000
	CLK = 1'b1;
    #10000; //3070000
	CLK = 1'b0;
    #10000; //3080000
	CLK = 1'b1;
    #10000; //3090000
	CLK = 1'b0;
    #10000; //3100000
	CLK = 1'b1;
    #10000; //3110000
	CLK = 1'b0;
    #10000; //3120000
	CLK = 1'b1;
    #10000; //3130000
	CLK = 1'b0;
    #10000; //3140000
	CLK = 1'b1;
    #10000; //3150000
	CLK = 1'b0;
    #10000; //3160000
	CLK = 1'b1;
    #10000; //3170000
	CLK = 1'b0;
    #10000; //3180000
	CLK = 1'b1;
    #10000; //3190000
	CLK = 1'b0;
    #10000; //3200000
	CLK = 1'b1;
    #10000; //3210000
	CLK = 1'b0;
    #10000; //3220000
	CLK = 1'b1;
    #10000; //3230000
	CLK = 1'b0;
    #10000; //3240000
	CLK = 1'b1;
    #10000; //3250000
	CLK = 1'b0;
    #10000; //3260000
	CLK = 1'b1;
    #10000; //3270000
	CLK = 1'b0;
    #10000; //3280000
	CLK = 1'b1;
    #10000; //3290000
	CLK = 1'b0;
    #10000; //3300000
	CLK = 1'b1;
    #10000; //3310000
	CLK = 1'b0;
    #10000; //3320000
	CLK = 1'b1;
    #10000; //3330000
	CLK = 1'b0;
    #10000; //3340000
	CLK = 1'b1;
    #10000; //3350000
	CLK = 1'b0;
    #10000; //3360000
	CLK = 1'b1;
    #10000; //3370000
	CLK = 1'b0;
    #10000; //3380000
	CLK = 1'b1;
    #10000; //3390000
	CLK = 1'b0;
    #10000; //3400000
	CLK = 1'b1;
    #10000; //3410000
	CLK = 1'b0;
    #10000; //3420000
	CLK = 1'b1;
    #10000; //3430000
	CLK = 1'b0;
    #10000; //3440000
	CLK = 1'b1;
    #10000; //3450000
	CLK = 1'b0;
    #10000; //3460000
	CLK = 1'b1;
    #10000; //3470000
	CLK = 1'b0;
    #10000; //3480000
	CLK = 1'b1;
    #10000; //3490000
	CLK = 1'b0;
    #10000; //3500000
	CLK = 1'b1;
    #10000; //3510000
	CLK = 1'b0;
    #10000; //3520000
	CLK = 1'b1;
    #10000; //3530000
	CLK = 1'b0;
    #10000; //3540000
	CLK = 1'b1;
    #10000; //3550000
	CLK = 1'b0;
    #10000; //3560000
	CLK = 1'b1;
    #10000; //3570000
	CLK = 1'b0;
    #10000; //3580000
	CLK = 1'b1;
    #10000; //3590000
	CLK = 1'b0;
    #10000; //3600000
	CLK = 1'b1;
    #10000; //3610000
	CLK = 1'b0;
    #10000; //3620000
	CLK = 1'b1;
    #10000; //3630000
	CLK = 1'b0;
    #10000; //3640000
	CLK = 1'b1;
    #10000; //3650000
	CLK = 1'b0;
    #10000; //3660000
	CLK = 1'b1;
    #10000; //3670000
	CLK = 1'b0;
    #10000; //3680000
	CLK = 1'b1;
    #10000; //3690000
	CLK = 1'b0;
    #10000; //3700000
	CLK = 1'b1;
    #10000; //3710000
	CLK = 1'b0;
    #10000; //3720000
	CLK = 1'b1;
    #10000; //3730000
	CLK = 1'b0;
    #10000; //3740000
	CLK = 1'b1;
    #10000; //3750000
	CLK = 1'b0;
    #10000; //3760000
	CLK = 1'b1;
    #10000; //3770000
	CLK = 1'b0;
    #10000; //3780000
	CLK = 1'b1;
    #10000; //3790000
	CLK = 1'b0;
    #10000; //3800000
	CLK = 1'b1;
    #10000; //3810000
	CLK = 1'b0;
    #10000; //3820000
	CLK = 1'b1;
    #10000; //3830000
	CLK = 1'b0;
    #10000; //3840000
	CLK = 1'b1;
    #10000; //3850000
	CLK = 1'b0;
    #10000; //3860000
	CLK = 1'b1;
    #10000; //3870000
	CLK = 1'b0;
    #10000; //3880000
	CLK = 1'b1;
    #10000; //3890000
	CLK = 1'b0;
    #10000; //3900000
	CLK = 1'b1;
    #10000; //3910000
	CLK = 1'b0;
    #10000; //3920000
	CLK = 1'b1;
    #10000; //3930000
	CLK = 1'b0;
    #10000; //3940000
	CLK = 1'b1;
    #10000; //3950000
	CLK = 1'b0;
    #10000; //3960000
	CLK = 1'b1;
    #10000; //3970000
	CLK = 1'b0;
    #10000; //3980000
	CLK = 1'b1;
    #10000; //3990000
	CLK = 1'b0;
    #10000; //4000000
	CLK = 1'b1;
    #10000; //4010000
	CLK = 1'b0;
    #10000; //4020000
	CLK = 1'b1;
    #10000; //4030000
	CLK = 1'b0;
    #10000; //4040000
	CLK = 1'b1;
    #10000; //4050000
	CLK = 1'b0;
    #10000; //4060000
	CLK = 1'b1;
    #10000; //4070000
	CLK = 1'b0;
    #10000; //4080000
	CLK = 1'b1;
    #10000; //4090000
	CLK = 1'b0;
    #10000; //4100000
	CLK = 1'b1;
    #10000; //4110000
	CLK = 1'b0;
    #10000; //4120000
	CLK = 1'b1;
    #10000; //4130000
	CLK = 1'b0;
    #10000; //4140000
	CLK = 1'b1;
    #10000; //4150000
	CLK = 1'b0;
    #10000; //4160000
	CLK = 1'b1;
    #10000; //4170000
	CLK = 1'b0;
    #10000; //4180000
	CLK = 1'b1;
    #10000; //4190000
	CLK = 1'b0;
    #10000; //4200000
	CLK = 1'b1;
    #10000; //4210000
	CLK = 1'b0;
    #10000; //4220000
	CLK = 1'b1;
    #10000; //4230000
	CLK = 1'b0;
    #10000; //4240000
	CLK = 1'b1;
    #10000; //4250000
	CLK = 1'b0;
    #10000; //4260000
	CLK = 1'b1;
    #10000; //4270000
	CLK = 1'b0;
    #10000; //4280000
	CLK = 1'b1;
    #10000; //4290000
	CLK = 1'b0;
    #10000; //4300000
	CLK = 1'b1;
    #10000; //4310000
	CLK = 1'b0;
    #10000; //4320000
	CLK = 1'b1;
    #10000; //4330000
	CLK = 1'b0;
    #10000; //4340000
	CLK = 1'b1;
    #10000; //4350000
	CLK = 1'b0;
    #10000; //4360000
	CLK = 1'b1;
    #10000; //4370000
	CLK = 1'b0;
    #10000; //4380000
	CLK = 1'b1;
    #10000; //4390000
	CLK = 1'b0;
    #10000; //4400000
	CLK = 1'b1;
    #10000; //4410000
	CLK = 1'b0;
    #10000; //4420000
	CLK = 1'b1;
    #10000; //4430000
	CLK = 1'b0;
    #10000; //4440000
	CLK = 1'b1;
    #10000; //4450000
	CLK = 1'b0;
    #10000; //4460000
	CLK = 1'b1;
    #10000; //4470000
	CLK = 1'b0;
    #10000; //4480000
	CLK = 1'b1;
    #10000; //4490000
	CLK = 1'b0;
    #10000; //4500000
	CLK = 1'b1;
    #10000; //4510000
	CLK = 1'b0;
    #10000; //4520000
	CLK = 1'b1;
    #10000; //4530000
	CLK = 1'b0;
    #10000; //4540000
	CLK = 1'b1;
    #10000; //4550000
	CLK = 1'b0;
    #10000; //4560000
	CLK = 1'b1;
    #10000; //4570000
	CLK = 1'b0;
    #10000; //4580000
	CLK = 1'b1;
    #10000; //4590000
	CLK = 1'b0;
    #10000; //4600000
	CLK = 1'b1;
    #10000; //4610000
	CLK = 1'b0;
    #10000; //4620000
	CLK = 1'b1;
    #10000; //4630000
	CLK = 1'b0;
    #10000; //4640000
	CLK = 1'b1;
    #10000; //4650000
	CLK = 1'b0;
    #10000; //4660000
	CLK = 1'b1;
    #10000; //4670000
	CLK = 1'b0;
    #10000; //4680000
	CLK = 1'b1;
    #10000; //4690000
	CLK = 1'b0;
    #10000; //4700000
	CLK = 1'b1;
    #10000; //4710000
	CLK = 1'b0;
    #10000; //4720000
	CLK = 1'b1;
    #10000; //4730000
	CLK = 1'b0;
    #10000; //4740000
	CLK = 1'b1;
    #10000; //4750000
	CLK = 1'b0;
    #10000; //4760000
	CLK = 1'b1;
    #10000; //4770000
	CLK = 1'b0;
    #10000; //4780000
	CLK = 1'b1;
    #10000; //4790000
	CLK = 1'b0;
    #10000; //4800000
	CLK = 1'b1;
    #10000; //4810000
	CLK = 1'b0;
    #10000; //4820000
	CLK = 1'b1;
    #10000; //4830000
	CLK = 1'b0;
    #10000; //4840000
	CLK = 1'b1;
    #10000; //4850000
	CLK = 1'b0;
    #10000; //4860000
	CLK = 1'b1;
    #10000; //4870000
	CLK = 1'b0;
    #10000; //4880000
	CLK = 1'b1;
    #10000; //4890000
	CLK = 1'b0;
    #10000; //4900000
	CLK = 1'b1;
    #10000; //4910000
	CLK = 1'b0;
    #10000; //4920000
	CLK = 1'b1;
    #10000; //4930000
	CLK = 1'b0;
    #10000; //4940000
	CLK = 1'b1;
    #10000; //4950000
	CLK = 1'b0;
    #10000; //4960000
	CLK = 1'b1;
    #10000; //4970000
	CLK = 1'b0;
    #10000; //4980000
	CLK = 1'b1;
    #10000; //4990000
	CLK = 1'b0;
    #10000; //5000000
	CLK = 1'b1;
    #10000; //5010000
	CLK = 1'b0;
    #10000; //5020000
	CLK = 1'b1;
    #10000; //5030000
	CLK = 1'b0;
    #10000; //5040000
	CLK = 1'b1;
    #10000; //5050000
	CLK = 1'b0;
    #10000; //5060000
	CLK = 1'b1;
    #10000; //5070000
	CLK = 1'b0;
    #10000; //5080000
	CLK = 1'b1;
    #10000; //5090000
	CLK = 1'b0;
    #10000; //5100000
	CLK = 1'b1;
    #10000; //5110000
	CLK = 1'b0;
    #10000; //5120000
	CLK = 1'b1;
    #10000; //5130000
	CLK = 1'b0;
    #10000; //5140000
	CLK = 1'b1;
    #10000; //5150000
	CLK = 1'b0;
    #10000; //5160000
	CLK = 1'b1;
    #10000; //5170000
	CLK = 1'b0;
    #10000; //5180000
	CLK = 1'b1;
    #10000; //5190000
	CLK = 1'b0;
    #10000; //5200000
	CLK = 1'b1;
    #10000; //5210000
	CLK = 1'b0;
    #10000; //5220000
	CLK = 1'b1;
    #10000; //5230000
	CLK = 1'b0;
    #10000; //5240000
	CLK = 1'b1;
    #10000; //5250000
	CLK = 1'b0;
    #10000; //5260000
	CLK = 1'b1;
    #10000; //5270000
	CLK = 1'b0;
    #10000; //5280000
	CLK = 1'b1;
    #10000; //5290000
	CLK = 1'b0;
    #10000; //5300000
	CLK = 1'b1;
    #10000; //5310000
	CLK = 1'b0;
    #10000; //5320000
	CLK = 1'b1;
    #10000; //5330000
	CLK = 1'b0;
    #10000; //5340000
	CLK = 1'b1;
    #10000; //5350000
	CLK = 1'b0;
    #10000; //5360000
	CLK = 1'b1;
    #10000; //5370000
	CLK = 1'b0;
    #10000; //5380000
	CLK = 1'b1;
    #10000; //5390000
	CLK = 1'b0;
    #10000; //5400000
	CLK = 1'b1;
    #10000; //5410000
	CLK = 1'b0;
    #10000; //5420000
	CLK = 1'b1;
    #10000; //5430000
	CLK = 1'b0;
    #10000; //5440000
	CLK = 1'b1;
    #10000; //5450000
	CLK = 1'b0;
    #10000; //5460000
	CLK = 1'b1;
    #10000; //5470000
	CLK = 1'b0;
    #10000; //5480000
	CLK = 1'b1;
    #10000; //5490000
	CLK = 1'b0;
    #10000; //5500000
	CLK = 1'b1;
    #10000; //5510000
	CLK = 1'b0;
    #10000; //5520000
	CLK = 1'b1;
    #10000; //5530000
	CLK = 1'b0;
    #10000; //5540000
	CLK = 1'b1;
    #10000; //5550000
	CLK = 1'b0;
    #10000; //5560000
	CLK = 1'b1;
    #10000; //5570000
	CLK = 1'b0;
    #10000; //5580000
	CLK = 1'b1;
    #10000; //5590000
	CLK = 1'b0;
    #10000; //5600000
	CLK = 1'b1;
    #10000; //5610000
	CLK = 1'b0;
    #10000; //5620000
	CLK = 1'b1;
    #10000; //5630000
	CLK = 1'b0;
    #10000; //5640000
	CLK = 1'b1;
    #10000; //5650000
	CLK = 1'b0;
    #10000; //5660000
	CLK = 1'b1;
    #10000; //5670000
	CLK = 1'b0;
    #10000; //5680000
	CLK = 1'b1;
    #10000; //5690000
	CLK = 1'b0;
    #10000; //5700000
	CLK = 1'b1;
    #10000; //5710000
	CLK = 1'b0;
    #10000; //5720000
	CLK = 1'b1;
    #10000; //5730000
	CLK = 1'b0;
    #10000; //5740000
	CLK = 1'b1;
    #10000; //5750000
	CLK = 1'b0;
    #10000; //5760000
	CLK = 1'b1;
    #10000; //5770000
	CLK = 1'b0;
    #10000; //5780000
	CLK = 1'b1;
    #10000; //5790000
	CLK = 1'b0;
    #10000; //5800000
	CLK = 1'b1;
    #10000; //5810000
	CLK = 1'b0;
    #10000; //5820000
	CLK = 1'b1;
    #10000; //5830000
	CLK = 1'b0;
    #10000; //5840000
	CLK = 1'b1;
    #10000; //5850000
	CLK = 1'b0;
    #10000; //5860000
	CLK = 1'b1;
    #10000; //5870000
	CLK = 1'b0;
    #10000; //5880000
	CLK = 1'b1;
    #10000; //5890000
	CLK = 1'b0;
    #10000; //5900000
	CLK = 1'b1;
    #10000; //5910000
	CLK = 1'b0;
    #10000; //5920000
	CLK = 1'b1;
    #10000; //5930000
	CLK = 1'b0;
    #10000; //5940000
	CLK = 1'b1;
    #10000; //5950000
	CLK = 1'b0;
    #10000; //5960000
	CLK = 1'b1;
    #10000; //5970000
	CLK = 1'b0;
    #10000; //5980000
	CLK = 1'b1;
    #10000; //5990000
	CLK = 1'b0;
    #10000; //6000000
	CLK = 1'b1;
    #10000; //6010000
	CLK = 1'b0;
    #10000; //6020000
	CLK = 1'b1;
    #10000; //6030000
	CLK = 1'b0;
    #10000; //6040000
	CLK = 1'b1;
    #10000; //6050000
	CLK = 1'b0;
    #10000; //6060000
	CLK = 1'b1;
    #10000; //6070000
	CLK = 1'b0;
    #10000; //6080000
	CLK = 1'b1;
    #10000; //6090000
	CLK = 1'b0;
    #10000; //6100000
	CLK = 1'b1;
    #10000; //6110000
	CLK = 1'b0;
    #10000; //6120000
	CLK = 1'b1;
    #10000; //6130000
	CLK = 1'b0;
    #10000; //6140000
	CLK = 1'b1;
    #10000; //6150000
	CLK = 1'b0;
    #10000; //6160000
	CLK = 1'b1;
    #10000; //6170000
	CLK = 1'b0;
    #10000; //6180000
	CLK = 1'b1;
    #10000; //6190000
	CLK = 1'b0;
    #10000; //6200000
	CLK = 1'b1;
    #10000; //6210000
	CLK = 1'b0;
    #10000; //6220000
	CLK = 1'b1;
    #10000; //6230000
	CLK = 1'b0;
    #10000; //6240000
	CLK = 1'b1;
    #10000; //6250000
	CLK = 1'b0;
    #10000; //6260000
	CLK = 1'b1;
    #10000; //6270000
	CLK = 1'b0;
    #10000; //6280000
	CLK = 1'b1;
    #10000; //6290000
	CLK = 1'b0;
    #10000; //6300000
	CLK = 1'b1;
    #10000; //6310000
	CLK = 1'b0;
    #10000; //6320000
	CLK = 1'b1;
    #10000; //6330000
	CLK = 1'b0;
    #10000; //6340000
	CLK = 1'b1;
    #10000; //6350000
	CLK = 1'b0;
    #10000; //6360000
	CLK = 1'b1;
    #10000; //6370000
	CLK = 1'b0;
    #10000; //6380000
	CLK = 1'b1;
    #10000; //6390000
	CLK = 1'b0;
    #10000; //6400000
	CLK = 1'b1;
    #10000; //6410000
	CLK = 1'b0;
    #10000; //6420000
	CLK = 1'b1;
    #10000; //6430000
	CLK = 1'b0;
    #10000; //6440000
	CLK = 1'b1;
    #10000; //6450000
	CLK = 1'b0;
    #10000; //6460000
	CLK = 1'b1;
    #10000; //6470000
	CLK = 1'b0;
    #10000; //6480000
	CLK = 1'b1;
    #10000; //6490000
	CLK = 1'b0;
    #10000; //6500000
	CLK = 1'b1;
    #10000; //6510000
	CLK = 1'b0;
    #10000; //6520000
	CLK = 1'b1;
    #10000; //6530000
	CLK = 1'b0;
    #10000; //6540000
	CLK = 1'b1;
    #10000; //6550000
	CLK = 1'b0;
    #10000; //6560000
	CLK = 1'b1;
    #10000; //6570000
	CLK = 1'b0;
    #10000; //6580000
	CLK = 1'b1;
    #10000; //6590000
	CLK = 1'b0;
    #10000; //6600000
	CLK = 1'b1;
    #10000; //6610000
	CLK = 1'b0;
    #10000; //6620000
	CLK = 1'b1;
    #10000; //6630000
	CLK = 1'b0;
    #10000; //6640000
	CLK = 1'b1;
    #10000; //6650000
	CLK = 1'b0;
    #10000; //6660000
	CLK = 1'b1;
    #10000; //6670000
	CLK = 1'b0;
    #10000; //6680000
	CLK = 1'b1;
    #10000; //6690000
	CLK = 1'b0;
    #10000; //6700000
	CLK = 1'b1;
    #10000; //6710000
	CLK = 1'b0;
    #10000; //6720000
	CLK = 1'b1;
    #10000; //6730000
	CLK = 1'b0;
    #10000; //6740000
	CLK = 1'b1;
    #10000; //6750000
	CLK = 1'b0;
    #10000; //6760000
	CLK = 1'b1;
    #10000; //6770000
	CLK = 1'b0;
    #10000; //6780000
	CLK = 1'b1;
    #10000; //6790000
	CLK = 1'b0;
    #10000; //6800000
	CLK = 1'b1;
    #10000; //6810000
	CLK = 1'b0;
    #10000; //6820000
	CLK = 1'b1;
    #10000; //6830000
	CLK = 1'b0;
    #10000; //6840000
	CLK = 1'b1;
    #10000; //6850000
	CLK = 1'b0;
    #10000; //6860000
	CLK = 1'b1;
    #10000; //6870000
	CLK = 1'b0;
    #10000; //6880000
	CLK = 1'b1;
    #10000; //6890000
	CLK = 1'b0;
    #10000; //6900000
	CLK = 1'b1;
    #10000; //6910000
	CLK = 1'b0;
    #10000; //6920000
	CLK = 1'b1;
    #10000; //6930000
	CLK = 1'b0;
    #10000; //6940000
	CLK = 1'b1;
    #10000; //6950000
	CLK = 1'b0;
    #10000; //6960000
	CLK = 1'b1;
    #10000; //6970000
	CLK = 1'b0;
    #10000; //6980000
	CLK = 1'b1;
    #10000; //6990000
	CLK = 1'b0;
    #10000; //7000000
	CLK = 1'b1;
    #10000; //7010000
	CLK = 1'b0;
    #10000; //7020000
	CLK = 1'b1;
    #10000; //7030000
	CLK = 1'b0;
    #10000; //7040000
	CLK = 1'b1;
    #10000; //7050000
	CLK = 1'b0;
    #10000; //7060000
	CLK = 1'b1;
    #10000; //7070000
	CLK = 1'b0;
    #10000; //7080000
	CLK = 1'b1;
    #10000; //7090000
	CLK = 1'b0;
    #10000; //7100000
	CLK = 1'b1;
    #10000; //7110000
	CLK = 1'b0;
    #10000; //7120000
	CLK = 1'b1;
    #10000; //7130000
	CLK = 1'b0;
    #10000; //7140000
	CLK = 1'b1;
    #10000; //7150000
	CLK = 1'b0;
    #10000; //7160000
	CLK = 1'b1;
    #10000; //7170000
	CLK = 1'b0;
    #10000; //7180000
	CLK = 1'b1;
    #10000; //7190000
	CLK = 1'b0;
    #10000; //7200000
	CLK = 1'b1;
    #10000; //7210000
	CLK = 1'b0;
    #10000; //7220000
	CLK = 1'b1;
    #10000; //7230000
	CLK = 1'b0;
    #10000; //7240000
	CLK = 1'b1;
    #10000; //7250000
	CLK = 1'b0;
    #10000; //7260000
	CLK = 1'b1;
    #10000; //7270000
	CLK = 1'b0;
    #10000; //7280000
	CLK = 1'b1;
    #10000; //7290000
	CLK = 1'b0;
    #10000; //7300000
	CLK = 1'b1;
    #10000; //7310000
	CLK = 1'b0;
    #10000; //7320000
	CLK = 1'b1;
    #10000; //7330000
	CLK = 1'b0;
    #10000; //7340000
	CLK = 1'b1;
    #10000; //7350000
	CLK = 1'b0;
    #10000; //7360000
	CLK = 1'b1;
    #10000; //7370000
	CLK = 1'b0;
    #10000; //7380000
	CLK = 1'b1;
    #10000; //7390000
	CLK = 1'b0;
    #10000; //7400000
	CLK = 1'b1;
    #10000; //7410000
	CLK = 1'b0;
    #10000; //7420000
	CLK = 1'b1;
    #10000; //7430000
	CLK = 1'b0;
    #10000; //7440000
	CLK = 1'b1;
    #10000; //7450000
	CLK = 1'b0;
    #10000; //7460000
	CLK = 1'b1;
    #10000; //7470000
	CLK = 1'b0;
    #10000; //7480000
	CLK = 1'b1;
    #10000; //7490000
	CLK = 1'b0;
    #10000; //7500000
	CLK = 1'b1;
    #10000; //7510000
	CLK = 1'b0;
    #10000; //7520000
	CLK = 1'b1;
    #10000; //7530000
	CLK = 1'b0;
    #10000; //7540000
	CLK = 1'b1;
    #10000; //7550000
	CLK = 1'b0;
    #10000; //7560000
	CLK = 1'b1;
    #10000; //7570000
	CLK = 1'b0;
    #10000; //7580000
	CLK = 1'b1;
    #10000; //7590000
	CLK = 1'b0;
    #10000; //7600000
	CLK = 1'b1;
    #10000; //7610000
	CLK = 1'b0;
    #10000; //7620000
	CLK = 1'b1;
    #10000; //7630000
	CLK = 1'b0;
    #10000; //7640000
	CLK = 1'b1;
    #10000; //7650000
	CLK = 1'b0;
    #10000; //7660000
	CLK = 1'b1;
    #10000; //7670000
	CLK = 1'b0;
    #10000; //7680000
	CLK = 1'b1;
    #10000; //7690000
	CLK = 1'b0;
    #10000; //7700000
	CLK = 1'b1;
    #10000; //7710000
	CLK = 1'b0;
    #10000; //7720000
	CLK = 1'b1;
    #10000; //7730000
	CLK = 1'b0;
    #10000; //7740000
	CLK = 1'b1;
    #10000; //7750000
	CLK = 1'b0;
    #10000; //7760000
	CLK = 1'b1;
    #10000; //7770000
	CLK = 1'b0;
    #10000; //7780000
	CLK = 1'b1;
    #10000; //7790000
	CLK = 1'b0;
    #10000; //7800000
	CLK = 1'b1;
    #10000; //7810000
	CLK = 1'b0;
    #10000; //7820000
	CLK = 1'b1;
    #10000; //7830000
	CLK = 1'b0;
    #10000; //7840000
	CLK = 1'b1;
    #10000; //7850000
	CLK = 1'b0;
    #10000; //7860000
	CLK = 1'b1;
    #10000; //7870000
	CLK = 1'b0;
    #10000; //7880000
	CLK = 1'b1;
    #10000; //7890000
	CLK = 1'b0;
    #10000; //7900000
	CLK = 1'b1;
    #10000; //7910000
	CLK = 1'b0;
    #10000; //7920000
	CLK = 1'b1;
    #10000; //7930000
	CLK = 1'b0;
    #10000; //7940000
	CLK = 1'b1;
    #10000; //7950000
	CLK = 1'b0;
    #10000; //7960000
	CLK = 1'b1;
    #10000; //7970000
	CLK = 1'b0;
    #10000; //7980000
	CLK = 1'b1;
    #10000; //7990000
	CLK = 1'b0;
    #10000; //8000000
	CLK = 1'b1;
    #10000; //8010000
	CLK = 1'b0;
    #10000; //8020000
	CLK = 1'b1;
    #10000; //8030000
	CLK = 1'b0;
    #10000; //8040000
	CLK = 1'b1;
    #10000; //8050000
	CLK = 1'b0;
    #10000; //8060000
	CLK = 1'b1;
    #10000; //8070000
	CLK = 1'b0;
    #10000; //8080000
	CLK = 1'b1;
    #10000; //8090000
	CLK = 1'b0;
    #10000; //8100000
	CLK = 1'b1;
    #10000; //8110000
	CLK = 1'b0;
    #10000; //8120000
	CLK = 1'b1;
    #10000; //8130000
	CLK = 1'b0;
    #10000; //8140000
	CLK = 1'b1;
    #10000; //8150000
	CLK = 1'b0;
    #10000; //8160000
	CLK = 1'b1;
    #10000; //8170000
	CLK = 1'b0;
    #10000; //8180000
	CLK = 1'b1;
    #10000; //8190000
	CLK = 1'b0;
    #10000; //8200000
	CLK = 1'b1;
    #10000; //8210000
	CLK = 1'b0;
    #10000; //8220000
	CLK = 1'b1;
    #10000; //8230000
	CLK = 1'b0;
    #10000; //8240000
	CLK = 1'b1;
    #10000; //8250000
	CLK = 1'b0;
    #10000; //8260000
	CLK = 1'b1;
    #10000; //8270000
	CLK = 1'b0;
    #10000; //8280000
	CLK = 1'b1;
    #10000; //8290000
	CLK = 1'b0;
    #10000; //8300000
	CLK = 1'b1;
    #10000; //8310000
	CLK = 1'b0;
    #10000; //8320000
	CLK = 1'b1;
    #10000; //8330000
	CLK = 1'b0;
    #10000; //8340000
	CLK = 1'b1;
    #10000; //8350000
	CLK = 1'b0;
    #10000; //8360000
	CLK = 1'b1;
    #10000; //8370000
	CLK = 1'b0;
    #10000; //8380000
	CLK = 1'b1;
    #10000; //8390000
	CLK = 1'b0;
    #10000; //8400000
	CLK = 1'b1;
    #10000; //8410000
	CLK = 1'b0;
    #10000; //8420000
	CLK = 1'b1;
    #10000; //8430000
	CLK = 1'b0;
    #10000; //8440000
	CLK = 1'b1;
    #10000; //8450000
	CLK = 1'b0;
    #10000; //8460000
	CLK = 1'b1;
    #10000; //8470000
	CLK = 1'b0;
    #10000; //8480000
	CLK = 1'b1;
    #10000; //8490000
	CLK = 1'b0;
    #10000; //8500000
	CLK = 1'b1;
    #10000; //8510000
	CLK = 1'b0;
    #10000; //8520000
	CLK = 1'b1;
    #10000; //8530000
	CLK = 1'b0;
    #10000; //8540000
	CLK = 1'b1;
    #10000; //8550000
	CLK = 1'b0;
    #10000; //8560000
	CLK = 1'b1;
    #10000; //8570000
	CLK = 1'b0;
    #10000; //8580000
	CLK = 1'b1;
    #10000; //8590000
	CLK = 1'b0;
    #10000; //8600000
	CLK = 1'b1;
    #10000; //8610000
	CLK = 1'b0;
    #10000; //8620000
	CLK = 1'b1;
    #10000; //8630000
	CLK = 1'b0;
    #10000; //8640000
	CLK = 1'b1;
    #10000; //8650000
	CLK = 1'b0;
    #10000; //8660000
	CLK = 1'b1;
    #10000; //8670000
	CLK = 1'b0;
    #10000; //8680000
	CLK = 1'b1;
    #10000; //8690000
	CLK = 1'b0;
    #10000; //8700000
	CLK = 1'b1;
    #10000; //8710000
	CLK = 1'b0;
    #10000; //8720000
	CLK = 1'b1;
    #10000; //8730000
	CLK = 1'b0;
    #10000; //8740000
	CLK = 1'b1;
    #10000; //8750000
	CLK = 1'b0;
    #10000; //8760000
	CLK = 1'b1;
    #10000; //8770000
	CLK = 1'b0;
    #10000; //8780000
	CLK = 1'b1;
    #10000; //8790000
	CLK = 1'b0;
    #10000; //8800000
	CLK = 1'b1;
    #10000; //8810000
	CLK = 1'b0;
    #10000; //8820000
	CLK = 1'b1;
    #10000; //8830000
	CLK = 1'b0;
    #10000; //8840000
	CLK = 1'b1;
    #10000; //8850000
	CLK = 1'b0;
    #10000; //8860000
	CLK = 1'b1;
    #10000; //8870000
	CLK = 1'b0;
    #10000; //8880000
	CLK = 1'b1;
    #10000; //8890000
	CLK = 1'b0;
    #10000; //8900000
	CLK = 1'b1;
    #10000; //8910000
	CLK = 1'b0;
    #10000; //8920000
	CLK = 1'b1;
    #10000; //8930000
	CLK = 1'b0;
    #10000; //8940000
	CLK = 1'b1;
    #10000; //8950000
	CLK = 1'b0;
    #10000; //8960000
	CLK = 1'b1;
    #10000; //8970000
	CLK = 1'b0;
    #10000; //8980000
	CLK = 1'b1;
    #10000; //8990000
	CLK = 1'b0;
    #10000; //9000000
	CLK = 1'b1;
    #10000; //9010000
	CLK = 1'b0;
    #10000; //9020000
	CLK = 1'b1;
    #10000; //9030000
	CLK = 1'b0;
    #10000; //9040000
	CLK = 1'b1;
    #10000; //9050000
	CLK = 1'b0;
    #10000; //9060000
	CLK = 1'b1;
    #10000; //9070000
	CLK = 1'b0;
    #10000; //9080000
	CLK = 1'b1;
    #10000; //9090000
	CLK = 1'b0;
    #10000; //9100000
	CLK = 1'b1;
    #10000; //9110000
	CLK = 1'b0;
    #10000; //9120000
	CLK = 1'b1;
    #10000; //9130000
	CLK = 1'b0;
    #10000; //9140000
	CLK = 1'b1;
    #10000; //9150000
	CLK = 1'b0;
    #10000; //9160000
	CLK = 1'b1;
    #10000; //9170000
	CLK = 1'b0;
    #10000; //9180000
	CLK = 1'b1;
    #10000; //9190000
	CLK = 1'b0;
    #10000; //9200000
	CLK = 1'b1;
    #10000; //9210000
	CLK = 1'b0;
    #10000; //9220000
	CLK = 1'b1;
    #10000; //9230000
	CLK = 1'b0;
    #10000; //9240000
	CLK = 1'b1;
    #10000; //9250000
	CLK = 1'b0;
    #10000; //9260000
	CLK = 1'b1;
    #10000; //9270000
	CLK = 1'b0;
    #10000; //9280000
	CLK = 1'b1;
    #10000; //9290000
	CLK = 1'b0;
    #10000; //9300000
	CLK = 1'b1;
    #10000; //9310000
	CLK = 1'b0;
    #10000; //9320000
	CLK = 1'b1;
    #10000; //9330000
	CLK = 1'b0;
    #5000; //9340000
	NI = 4'b0001;
    #5000; //9345000
	CLK = 1'b1;
    #10000; //9350000
	CLK = 1'b0;
    #10000; //9360000
	CLK = 1'b1;
    #10000; //9370000
	CLK = 1'b0;
    #10000; //9380000
	CLK = 1'b1;
    #10000; //9390000
	CLK = 1'b0;
    #10000; //9400000
	CLK = 1'b1;
    #10000; //9410000
	CLK = 1'b0;
    #10000; //9420000
	CLK = 1'b1;
    #10000; //9430000
	CLK = 1'b0;
    #10000; //9440000
	CLK = 1'b1;
    #10000; //9450000
	CLK = 1'b0;
    #10000; //9460000
	CLK = 1'b1;
    #10000; //9470000
	CLK = 1'b0;
    #10000; //9480000
	CLK = 1'b1;
    #10000; //9490000
	CLK = 1'b0;
    #10000; //9500000
	CLK = 1'b1;
    #10000; //9510000
	CLK = 1'b0;
    #10000; //9520000
	CLK = 1'b1;
    #10000; //9530000
	CLK = 1'b0;
    #10000; //9540000
	CLK = 1'b1;
    #10000; //9550000
	CLK = 1'b0;
    #10000; //9560000
	CLK = 1'b1;
    #10000; //9570000
	CLK = 1'b0;
    #10000; //9580000
	CLK = 1'b1;
    #10000; //9590000
	CLK = 1'b0;
    #10000; //9600000
	CLK = 1'b1;
    #10000; //9610000
	CLK = 1'b0;
    #10000; //9620000
	CLK = 1'b1;
    #10000; //9630000
	CLK = 1'b0;
    #10000; //9640000
	CLK = 1'b1;
    #10000; //9650000
	CLK = 1'b0;
    #10000; //9660000
	CLK = 1'b1;
    #10000; //9670000
	CLK = 1'b0;
    #10000; //9680000
	CLK = 1'b1;
    #10000; //9690000
	CLK = 1'b0;
    #10000; //9700000
	CLK = 1'b1;
    #10000; //9710000
	CLK = 1'b0;
    #10000; //9720000
	CLK = 1'b1;
    #10000; //9730000
	CLK = 1'b0;
    #10000; //9740000
	CLK = 1'b1;
    #10000; //9750000
	CLK = 1'b0;
    #10000; //9760000
	CLK = 1'b1;
    #10000; //9770000
	CLK = 1'b0;
    #10000; //9780000
	CLK = 1'b1;
    #10000; //9790000
	CLK = 1'b0;
    #10000; //9800000
	CLK = 1'b1;
    #10000; //9810000
	CLK = 1'b0;
    #10000; //9820000
	CLK = 1'b1;
    #10000; //9830000
	CLK = 1'b0;
    #10000; //9840000
	CLK = 1'b1;
    #10000; //9850000
	CLK = 1'b0;
    #10000; //9860000
	CLK = 1'b1;
    #10000; //9870000
	CLK = 1'b0;
    #10000; //9880000
	CLK = 1'b1;
    #10000; //9890000
	CLK = 1'b0;
    #10000; //9900000
	CLK = 1'b1;
    #10000; //9910000
	CLK = 1'b0;
    #10000; //9920000
	CLK = 1'b1;
    #10000; //9930000
	CLK = 1'b0;
    #10000; //9940000
	CLK = 1'b1;
    #10000; //9950000
	CLK = 1'b0;
    #10000; //9960000
	CLK = 1'b1;
    #10000; //9970000
	CLK = 1'b0;
    #10000; //9980000
	CLK = 1'b1;
    #10000; //9990000
	CLK = 1'b0;
    #10000; //10000000
	CLK = 1'b1;
    #10000; //10010000
	CLK = 1'b0;
    #10000; //10020000
	CLK = 1'b1;
    #10000; //10030000
	CLK = 1'b0;
    #10000; //10040000
	CLK = 1'b1;
    #10000; //10050000
	CLK = 1'b0;
    #10000; //10060000
	CLK = 1'b1;
    #10000; //10070000
	CLK = 1'b0;
    #10000; //10080000
	CLK = 1'b1;
    #10000; //10090000
	CLK = 1'b0;
    #10000; //10100000
	CLK = 1'b1;
    #10000; //10110000
	CLK = 1'b0;
    #10000; //10120000
	CLK = 1'b1;
    #10000; //10130000
	CLK = 1'b0;
    #10000; //10140000
	CLK = 1'b1;
    #10000; //10150000
	CLK = 1'b0;
    #10000; //10160000
	CLK = 1'b1;
    #10000; //10170000
	CLK = 1'b0;
    #10000; //10180000
	CLK = 1'b1;
    #10000; //10190000
	CLK = 1'b0;
    #10000; //10200000
	CLK = 1'b1;
    #10000; //10210000
	CLK = 1'b0;
    #10000; //10220000
	CLK = 1'b1;
    #10000; //10230000
	CLK = 1'b0;
    #10000; //10240000
	CLK = 1'b1;
    #10000; //10250000
	CLK = 1'b0;
    #10000; //10260000
	CLK = 1'b1;
    #10000; //10270000
	CLK = 1'b0;
    #10000; //10280000
	CLK = 1'b1;
    #10000; //10290000
	CLK = 1'b0;
    #10000; //10300000
	CLK = 1'b1;
    #10000; //10310000
	CLK = 1'b0;
    #10000; //10320000
	CLK = 1'b1;
    #10000; //10330000
	CLK = 1'b0;
    #10000; //10340000
	CLK = 1'b1;
    #10000; //10350000
	CLK = 1'b0;
    #10000; //10360000
	CLK = 1'b1;
    #10000; //10370000
	CLK = 1'b0;
    #10000; //10380000
	CLK = 1'b1;
    #10000; //10390000
	CLK = 1'b0;
    #10000; //10400000
	CLK = 1'b1;
    #10000; //10410000
	CLK = 1'b0;
    #10000; //10420000
	CLK = 1'b1;
    #10000; //10430000
	CLK = 1'b0;
    #10000; //10440000
	CLK = 1'b1;
    #10000; //10450000
	CLK = 1'b0;
    #10000; //10460000
	CLK = 1'b1;
    #10000; //10470000
	CLK = 1'b0;
    #10000; //10480000
	CLK = 1'b1;
    #10000; //10490000
	CLK = 1'b0;
    #10000; //10500000
	CLK = 1'b1;
    #10000; //10510000
	CLK = 1'b0;
    #10000; //10520000
	CLK = 1'b1;
    #10000; //10530000
	CLK = 1'b0;
    #10000; //10540000
	CLK = 1'b1;
    #10000; //10550000
	CLK = 1'b0;
    #10000; //10560000
	CLK = 1'b1;
    #10000; //10570000
	CLK = 1'b0;
    #10000; //10580000
	CLK = 1'b1;
    #10000; //10590000
	CLK = 1'b0;
    #10000; //10600000
	CLK = 1'b1;
    #10000; //10610000
	CLK = 1'b0;
    #10000; //10620000
	CLK = 1'b1;
    #10000; //10630000
	CLK = 1'b0;
    #10000; //10640000
	CLK = 1'b1;
    #10000; //10650000
	CLK = 1'b0;
    #10000; //10660000
	CLK = 1'b1;
    #10000; //10670000
	CLK = 1'b0;
    #10000; //10680000
	CLK = 1'b1;
    #10000; //10690000
	CLK = 1'b0;
    #10000; //10700000
	CLK = 1'b1;
    #10000; //10710000
	CLK = 1'b0;
    #10000; //10720000
	CLK = 1'b1;
    #10000; //10730000
	CLK = 1'b0;
    #10000; //10740000
	CLK = 1'b1;
    #10000; //10750000
	CLK = 1'b0;
    #10000; //10760000
	CLK = 1'b1;
    #10000; //10770000
	CLK = 1'b0;
    #10000; //10780000
	CLK = 1'b1;
    #10000; //10790000
	CLK = 1'b0;
    #10000; //10800000
	CLK = 1'b1;
    #10000; //10810000
	CLK = 1'b0;
    #10000; //10820000
	CLK = 1'b1;
    #10000; //10830000
	CLK = 1'b0;
    #10000; //10840000
	CLK = 1'b1;
    #10000; //10850000
	CLK = 1'b0;
    #10000; //10860000
	CLK = 1'b1;
    #10000; //10870000
	CLK = 1'b0;
    #10000; //10880000
	CLK = 1'b1;
    #10000; //10890000
	CLK = 1'b0;
    #10000; //10900000
	CLK = 1'b1;
    #10000; //10910000
	CLK = 1'b0;
    #10000; //10920000
	CLK = 1'b1;
    #10000; //10930000
	CLK = 1'b0;
    #10000; //10940000
	CLK = 1'b1;
    #10000; //10950000
	CLK = 1'b0;
    #10000; //10960000
	CLK = 1'b1;
    #10000; //10970000
	CLK = 1'b0;
    #10000; //10980000
	CLK = 1'b1;
    #10000; //10990000
	CLK = 1'b0;
    #10000; //11000000
	CLK = 1'b1;
    #10000; //11010000
	CLK = 1'b0;
    #10000; //11020000
	CLK = 1'b1;
    #10000; //11030000
	CLK = 1'b0;
    #10000; //11040000
	CLK = 1'b1;
    #10000; //11050000
	CLK = 1'b0;
    #10000; //11060000
	CLK = 1'b1;
    #10000; //11070000
	CLK = 1'b0;
    #10000; //11080000
	CLK = 1'b1;
    #10000; //11090000
	CLK = 1'b0;
    #10000; //11100000
	CLK = 1'b1;
    #10000; //11110000
	CLK = 1'b0;
    #10000; //11120000
	CLK = 1'b1;
    #10000; //11130000
	CLK = 1'b0;
    #10000; //11140000
	CLK = 1'b1;
    #10000; //11150000
	CLK = 1'b0;
    #10000; //11160000
	CLK = 1'b1;
    #10000; //11170000
	CLK = 1'b0;
    #10000; //11180000
	CLK = 1'b1;
    #10000; //11190000
	CLK = 1'b0;
    #10000; //11200000
	CLK = 1'b1;
    #10000; //11210000
	CLK = 1'b0;
    #10000; //11220000
	CLK = 1'b1;
    #10000; //11230000
	CLK = 1'b0;
    #10000; //11240000
	CLK = 1'b1;
    #10000; //11250000
	CLK = 1'b0;
    #10000; //11260000
	CLK = 1'b1;
    #10000; //11270000
	CLK = 1'b0;
    #10000; //11280000
	CLK = 1'b1;
    #10000; //11290000
	CLK = 1'b0;
    #10000; //11300000
	CLK = 1'b1;
    #10000; //11310000
	CLK = 1'b0;
    #10000; //11320000
	CLK = 1'b1;
    #10000; //11330000
	CLK = 1'b0;
    #10000; //11340000
	CLK = 1'b1;
    #10000; //11350000
	CLK = 1'b0;
    #10000; //11360000
	CLK = 1'b1;
    #10000; //11370000
	CLK = 1'b0;
    #10000; //11380000
	CLK = 1'b1;
    #10000; //11390000
	CLK = 1'b0;
    #10000; //11400000
	CLK = 1'b1;
    #10000; //11410000
	CLK = 1'b0;
    #10000; //11420000
	CLK = 1'b1;
    #10000; //11430000
	CLK = 1'b0;
    #10000; //11440000
	CLK = 1'b1;
    #10000; //11450000
	CLK = 1'b0;
    #10000; //11460000
	CLK = 1'b1;
    #10000; //11470000
	CLK = 1'b0;
    #10000; //11480000
	CLK = 1'b1;
    #10000; //11490000
	CLK = 1'b0;
    #10000; //11500000
	CLK = 1'b1;
    #10000; //11510000
	CLK = 1'b0;
    #10000; //11520000
	CLK = 1'b1;
    #10000; //11530000
	CLK = 1'b0;
    #10000; //11540000
	CLK = 1'b1;
    #10000; //11550000
	CLK = 1'b0;
    #10000; //11560000
	CLK = 1'b1;
    #10000; //11570000
	CLK = 1'b0;
    #10000; //11580000
	CLK = 1'b1;
    #10000; //11590000
	CLK = 1'b0;
    #10000; //11600000
	CLK = 1'b1;
    #10000; //11610000
	CLK = 1'b0;
    #10000; //11620000
	CLK = 1'b1;
    #10000; //11630000
	CLK = 1'b0;
    #10000; //11640000
	CLK = 1'b1;
    #10000; //11650000
	CLK = 1'b0;
    #10000; //11660000
	CLK = 1'b1;
    #10000; //11670000
	CLK = 1'b0;
    #10000; //11680000
	CLK = 1'b1;
    #10000; //11690000
	CLK = 1'b0;
    #10000; //11700000
	CLK = 1'b1;
    #10000; //11710000
	CLK = 1'b0;
    #10000; //11720000
	CLK = 1'b1;
    #10000; //11730000
	CLK = 1'b0;
    #10000; //11740000
	CLK = 1'b1;
    #10000; //11750000
	CLK = 1'b0;
    #10000; //11760000
	CLK = 1'b1;
    #10000; //11770000
	CLK = 1'b0;
    #10000; //11780000
	CLK = 1'b1;
    #10000; //11790000
	CLK = 1'b0;
    #10000; //11800000
	CLK = 1'b1;
    #10000; //11810000
	CLK = 1'b0;
    #10000; //11820000
	CLK = 1'b1;
    #10000; //11830000
	CLK = 1'b0;
    #10000; //11840000
	CLK = 1'b1;
    #10000; //11850000
	CLK = 1'b0;
    #10000; //11860000
	CLK = 1'b1;
    #10000; //11870000
	CLK = 1'b0;
    #10000; //11880000
	CLK = 1'b1;
    #10000; //11890000
	CLK = 1'b0;
    #10000; //11900000
	CLK = 1'b1;
    #10000; //11910000
	CLK = 1'b0;
    #10000; //11920000
	CLK = 1'b1;
    #10000; //11930000
	CLK = 1'b0;
    #10000; //11940000
	CLK = 1'b1;
    #10000; //11950000
	CLK = 1'b0;
    #10000; //11960000
	CLK = 1'b1;
    #10000; //11970000
	CLK = 1'b0;
    #10000; //11980000
	CLK = 1'b1;
    #10000; //11990000
	CLK = 1'b0;
    #10000; //12000000
	CLK = 1'b1;
    #10000; //12010000
	CLK = 1'b0;
    #10000; //12020000
	CLK = 1'b1;
    #10000; //12030000
	CLK = 1'b0;
    #10000; //12040000
	CLK = 1'b1;
    #10000; //12050000
	CLK = 1'b0;
    #10000; //12060000
	CLK = 1'b1;
    #10000; //12070000
	CLK = 1'b0;
    #10000; //12080000
	CLK = 1'b1;
    #10000; //12090000
	CLK = 1'b0;
    #10000; //12100000
	CLK = 1'b1;
    #10000; //12110000
	CLK = 1'b0;
    #10000; //12120000
	CLK = 1'b1;
    #10000; //12130000
	CLK = 1'b0;
    #10000; //12140000
	CLK = 1'b1;
    #10000; //12150000
	CLK = 1'b0;
    #10000; //12160000
	CLK = 1'b1;
    #10000; //12170000
	CLK = 1'b0;
    #10000; //12180000
	CLK = 1'b1;
    #10000; //12190000
	CLK = 1'b0;
    #10000; //12200000
	CLK = 1'b1;
    #10000; //12210000
	CLK = 1'b0;
    #10000; //12220000
	CLK = 1'b1;
    #10000; //12230000
	CLK = 1'b0;
    #10000; //12240000
	CLK = 1'b1;
    #10000; //12250000
	CLK = 1'b0;
    #10000; //12260000
	CLK = 1'b1;
    #10000; //12270000
	CLK = 1'b0;
    #10000; //12280000
	CLK = 1'b1;
    #10000; //12290000
	CLK = 1'b0;
    #10000; //12300000
	CLK = 1'b1;
    #10000; //12310000
	CLK = 1'b0;
    #10000; //12320000
	CLK = 1'b1;
    #10000; //12330000
	CLK = 1'b0;
    #10000; //12340000
	CLK = 1'b1;
    #10000; //12350000
	CLK = 1'b0;
    #10000; //12360000
	CLK = 1'b1;
    #10000; //12370000
	CLK = 1'b0;
    #10000; //12380000
	CLK = 1'b1;
    #10000; //12390000
	CLK = 1'b0;
    #10000; //12400000
	CLK = 1'b1;
    #10000; //12410000
	CLK = 1'b0;
    #10000; //12420000
	CLK = 1'b1;
    #10000; //12430000
	CLK = 1'b0;
    #10000; //12440000
	CLK = 1'b1;
    #10000; //12450000
	CLK = 1'b0;
    #10000; //12460000
	CLK = 1'b1;
    #10000; //12470000
	CLK = 1'b0;
    #10000; //12480000
	CLK = 1'b1;
    #10000; //12490000
	CLK = 1'b0;
    #10000; //12500000
	CLK = 1'b1;
    #10000; //12510000
	CLK = 1'b0;
    #10000; //12520000
	CLK = 1'b1;
    #10000; //12530000
	CLK = 1'b0;
    #10000; //12540000
	CLK = 1'b1;
    #10000; //12550000
	CLK = 1'b0;
    #10000; //12560000
	CLK = 1'b1;
    #10000; //12570000
	CLK = 1'b0;
    #10000; //12580000
	CLK = 1'b1;
    #10000; //12590000
	CLK = 1'b0;
    #10000; //12600000
	CLK = 1'b1;
    #10000; //12610000
	CLK = 1'b0;
    #10000; //12620000
	CLK = 1'b1;
    #10000; //12630000
	CLK = 1'b0;
    #10000; //12640000
	CLK = 1'b1;
    #10000; //12650000
	CLK = 1'b0;
    #10000; //12660000
	CLK = 1'b1;
    #10000; //12670000
	CLK = 1'b0;
    #10000; //12680000
	CLK = 1'b1;
    #10000; //12690000
	CLK = 1'b0;
    #10000; //12700000
	CLK = 1'b1;
    #10000; //12710000
	CLK = 1'b0;
    #10000; //12720000
	CLK = 1'b1;
    #10000; //12730000
	CLK = 1'b0;
    #10000; //12740000
	CLK = 1'b1;
    #10000; //12750000
	CLK = 1'b0;
    #10000; //12760000
	CLK = 1'b1;
    #10000; //12770000
	CLK = 1'b0;
    #10000; //12780000
	CLK = 1'b1;
    #10000; //12790000
	CLK = 1'b0;
    #10000; //12800000
	CLK = 1'b1;
    #10000; //12810000
	CLK = 1'b0;
    #10000; //12820000
	CLK = 1'b1;
    #10000; //12830000
	CLK = 1'b0;
    #10000; //12840000
	CLK = 1'b1;
    #10000; //12850000
	CLK = 1'b0;
    #10000; //12860000
	CLK = 1'b1;
    #10000; //12870000
	CLK = 1'b0;
    #10000; //12880000
	CLK = 1'b1;
    #10000; //12890000
	CLK = 1'b0;
    #10000; //12900000
	CLK = 1'b1;
    #10000; //12910000
	CLK = 1'b0;
    #10000; //12920000
	CLK = 1'b1;
    #10000; //12930000
	CLK = 1'b0;
    #10000; //12940000
	CLK = 1'b1;
    #10000; //12950000
	CLK = 1'b0;
    #10000; //12960000
	CLK = 1'b1;
    #10000; //12970000
	CLK = 1'b0;
    #10000; //12980000
	CLK = 1'b1;
    #10000; //12990000
	CLK = 1'b0;
    #10000; //13000000
	CLK = 1'b1;
    #10000; //13010000
	CLK = 1'b0;
    #10000; //13020000
	CLK = 1'b1;
    #10000; //13030000
	CLK = 1'b0;
    #10000; //13040000
	CLK = 1'b1;
    #10000; //13050000
	CLK = 1'b0;
    #10000; //13060000
	CLK = 1'b1;
    #10000; //13070000
	CLK = 1'b0;
    #10000; //13080000
	CLK = 1'b1;
    #10000; //13090000
	CLK = 1'b0;
    #10000; //13100000
	CLK = 1'b1;
    #10000; //13110000
	CLK = 1'b0;
    #10000; //13120000
	CLK = 1'b1;
    #10000; //13130000
	CLK = 1'b0;
    #10000; //13140000
	CLK = 1'b1;
    #10000; //13150000
	CLK = 1'b0;
    #10000; //13160000
	CLK = 1'b1;
    #10000; //13170000
	CLK = 1'b0;
    #10000; //13180000
	CLK = 1'b1;
    #10000; //13190000
	CLK = 1'b0;
    #10000; //13200000
	CLK = 1'b1;
    #10000; //13210000
	CLK = 1'b0;
    #10000; //13220000
	CLK = 1'b1;
    #10000; //13230000
	CLK = 1'b0;
    #10000; //13240000
	CLK = 1'b1;
    #10000; //13250000
	CLK = 1'b0;
    #10000; //13260000
	CLK = 1'b1;
    #10000; //13270000
	CLK = 1'b0;
    #10000; //13280000
	CLK = 1'b1;
    #10000; //13290000
	CLK = 1'b0;
    #10000; //13300000
	CLK = 1'b1;
    #10000; //13310000
	CLK = 1'b0;
    #10000; //13320000
	CLK = 1'b1;
    #10000; //13330000
	CLK = 1'b0;
    #10000; //13340000
	CLK = 1'b1;
    #10000; //13350000
	CLK = 1'b0;
    #10000; //13360000
	CLK = 1'b1;
    #10000; //13370000
	CLK = 1'b0;
    #10000; //13380000
	CLK = 1'b1;
    #10000; //13390000
	CLK = 1'b0;
    #10000; //13400000
	CLK = 1'b1;
    #10000; //13410000
	CLK = 1'b0;
    #10000; //13420000
	CLK = 1'b1;
    #10000; //13430000
	CLK = 1'b0;
    #10000; //13440000
	CLK = 1'b1;
    #10000; //13450000
	CLK = 1'b0;
    #10000; //13460000
	CLK = 1'b1;
    #10000; //13470000
	CLK = 1'b0;
    #10000; //13480000
	CLK = 1'b1;
    #10000; //13490000
	CLK = 1'b0;
    #10000; //13500000
	CLK = 1'b1;
    #10000; //13510000
	CLK = 1'b0;
    #10000; //13520000
	CLK = 1'b1;
    #10000; //13530000
	CLK = 1'b0;
    #10000; //13540000
	CLK = 1'b1;
    #10000; //13550000
	CLK = 1'b0;
    #10000; //13560000
	CLK = 1'b1;
    #10000; //13570000
	CLK = 1'b0;
    #10000; //13580000
	CLK = 1'b1;
    #10000; //13590000
	CLK = 1'b0;
    #10000; //13600000
	CLK = 1'b1;
    #10000; //13610000
	CLK = 1'b0;
    #10000; //13620000
	CLK = 1'b1;
    #10000; //13630000
	CLK = 1'b0;
    #10000; //13640000
	CLK = 1'b1;
    #10000; //13650000
	CLK = 1'b0;
    #10000; //13660000
	CLK = 1'b1;
    #10000; //13670000
	CLK = 1'b0;
    #10000; //13680000
	CLK = 1'b1;
    #10000; //13690000
	CLK = 1'b0;
    #10000; //13700000
	CLK = 1'b1;
    #10000; //13710000
	CLK = 1'b0;
    #10000; //13720000
	CLK = 1'b1;
    #10000; //13730000
	CLK = 1'b0;
    #10000; //13740000
	CLK = 1'b1;
    #10000; //13750000
	CLK = 1'b0;
    #10000; //13760000
	CLK = 1'b1;
    #10000; //13770000
	CLK = 1'b0;
    #10000; //13780000
	CLK = 1'b1;
    #10000; //13790000
	CLK = 1'b0;
    #10000; //13800000
	CLK = 1'b1;
    #10000; //13810000
	CLK = 1'b0;
    #10000; //13820000
	CLK = 1'b1;
    #10000; //13830000
	CLK = 1'b0;
    #10000; //13840000
	CLK = 1'b1;
    #10000; //13850000
	CLK = 1'b0;
    #10000; //13860000
	CLK = 1'b1;
    #10000; //13870000
	CLK = 1'b0;
    #10000; //13880000
	CLK = 1'b1;
    #10000; //13890000
	CLK = 1'b0;
    #10000; //13900000
	CLK = 1'b1;
    #10000; //13910000
	CLK = 1'b0;
    #10000; //13920000
	CLK = 1'b1;
    #10000; //13930000
	CLK = 1'b0;
    #10000; //13940000
	CLK = 1'b1;
    #10000; //13950000
	CLK = 1'b0;
    #10000; //13960000
	CLK = 1'b1;
    #10000; //13970000
	CLK = 1'b0;
    #10000; //13980000
	CLK = 1'b1;
    #10000; //13990000
	CLK = 1'b0;
    #10000; //14000000
	CLK = 1'b1;
    #10000; //14010000
	CLK = 1'b0;
    #10000; //14020000
	CLK = 1'b1;
    #10000; //14030000
	CLK = 1'b0;
    #10000; //14040000
	CLK = 1'b1;
    #10000; //14050000
	CLK = 1'b0;
    #10000; //14060000
	CLK = 1'b1;
    #10000; //14070000
	CLK = 1'b0;
    #10000; //14080000
	CLK = 1'b1;
    #10000; //14090000
	CLK = 1'b0;
    #10000; //14100000
	CLK = 1'b1;
    #10000; //14110000
	CLK = 1'b0;
    #10000; //14120000
	CLK = 1'b1;
    #10000; //14130000
	CLK = 1'b0;
    #10000; //14140000
	CLK = 1'b1;
    #10000; //14150000
	CLK = 1'b0;
    #10000; //14160000
	CLK = 1'b1;
    #10000; //14170000
	CLK = 1'b0;
    #10000; //14180000
	CLK = 1'b1;
    #10000; //14190000
	CLK = 1'b0;
    #10000; //14200000
	CLK = 1'b1;
    #10000; //14210000
	CLK = 1'b0;
    #10000; //14220000
	CLK = 1'b1;
    #10000; //14230000
	CLK = 1'b0;
    #10000; //14240000
	CLK = 1'b1;
    #10000; //14250000
	CLK = 1'b0;
    #10000; //14260000
	CLK = 1'b1;
    #10000; //14270000
	CLK = 1'b0;
    #10000; //14280000
	CLK = 1'b1;
    #10000; //14290000
	CLK = 1'b0;
    #10000; //14300000
	CLK = 1'b1;
    #10000; //14310000
	CLK = 1'b0;
    #10000; //14320000
	CLK = 1'b1;
    #10000; //14330000
	CLK = 1'b0;
    #10000; //14340000
	CLK = 1'b1;
    #10000; //14350000
	CLK = 1'b0;
    #10000; //14360000
	CLK = 1'b1;
    #10000; //14370000
	CLK = 1'b0;
    #10000; //14380000
	CLK = 1'b1;
    #10000; //14390000
	CLK = 1'b0;
    #10000; //14400000
	CLK = 1'b1;
    #10000; //14410000
	CLK = 1'b0;
    #10000; //14420000
	CLK = 1'b1;
    #10000; //14430000
	CLK = 1'b0;
    #10000; //14440000
	CLK = 1'b1;
    #10000; //14450000
	CLK = 1'b0;
    #10000; //14460000
	CLK = 1'b1;
    #10000; //14470000
	CLK = 1'b0;
    #10000; //14480000
	CLK = 1'b1;
    #10000; //14490000
	CLK = 1'b0;
    #10000; //14500000
	CLK = 1'b1;
    #10000; //14510000
	CLK = 1'b0;
    #10000; //14520000
	CLK = 1'b1;
    #10000; //14530000
	CLK = 1'b0;
    #10000; //14540000
	CLK = 1'b1;
    #10000; //14550000
	CLK = 1'b0;
    #10000; //14560000
	CLK = 1'b1;
    #10000; //14570000
	CLK = 1'b0;
    #10000; //14580000
	CLK = 1'b1;
    #10000; //14590000
	CLK = 1'b0;
    #10000; //14600000
	CLK = 1'b1;
    #10000; //14610000
	CLK = 1'b0;
    #10000; //14620000
	CLK = 1'b1;
    #10000; //14630000
	CLK = 1'b0;
    #10000; //14640000
	CLK = 1'b1;
    #10000; //14650000
	CLK = 1'b0;
    #10000; //14660000
	CLK = 1'b1;
    #10000; //14670000
	CLK = 1'b0;
    #10000; //14680000
	CLK = 1'b1;
    #10000; //14690000
	CLK = 1'b0;
    #10000; //14700000
	CLK = 1'b1;
    #10000; //14710000
	CLK = 1'b0;
    #10000; //14720000
	CLK = 1'b1;
    #10000; //14730000
	CLK = 1'b0;
    #10000; //14740000
	CLK = 1'b1;
    #10000; //14750000
	CLK = 1'b0;
    #10000; //14760000
	CLK = 1'b1;
    #10000; //14770000
	CLK = 1'b0;
    #10000; //14780000
	CLK = 1'b1;
    #10000; //14790000
	CLK = 1'b0;
    #10000; //14800000
	CLK = 1'b1;
    #10000; //14810000
	CLK = 1'b0;
    #10000; //14820000
	CLK = 1'b1;
    #10000; //14830000
	CLK = 1'b0;
    #10000; //14840000
	CLK = 1'b1;
    #10000; //14850000
	CLK = 1'b0;
    #10000; //14860000
	CLK = 1'b1;
    #10000; //14870000
	CLK = 1'b0;
    #10000; //14880000
	CLK = 1'b1;
    #10000; //14890000
	CLK = 1'b0;
    #10000; //14900000
	CLK = 1'b1;
    #10000; //14910000
	CLK = 1'b0;
    #10000; //14920000
	CLK = 1'b1;
    #10000; //14930000
	CLK = 1'b0;
    #10000; //14940000
	CLK = 1'b1;
    #10000; //14950000
	CLK = 1'b0;
    #10000; //14960000
	CLK = 1'b1;
    #10000; //14970000
	CLK = 1'b0;
    #10000; //14980000
	CLK = 1'b1;
    #10000; //14990000
	CLK = 1'b0;
    #10000; //15000000
	CLK = 1'b1;
    #10000; //15010000
	CLK = 1'b0;
    #10000; //15020000
	CLK = 1'b1;
    #10000; //15030000
	CLK = 1'b0;
    #10000; //15040000
	CLK = 1'b1;
    #10000; //15050000
	CLK = 1'b0;
    #10000; //15060000
	CLK = 1'b1;
    #10000; //15070000
	CLK = 1'b0;
    #10000; //15080000
	CLK = 1'b1;
    #10000; //15090000
	CLK = 1'b0;
    #10000; //15100000
	CLK = 1'b1;
    #10000; //15110000
	CLK = 1'b0;
    #10000; //15120000
	CLK = 1'b1;
    #10000; //15130000
	CLK = 1'b0;
    #10000; //15140000
	CLK = 1'b1;
    #10000; //15150000
	CLK = 1'b0;
    #10000; //15160000
	CLK = 1'b1;
    #10000; //15170000
	CLK = 1'b0;
    #10000; //15180000
	CLK = 1'b1;
    #10000; //15190000
	CLK = 1'b0;
    #10000; //15200000
	CLK = 1'b1;
    #10000; //15210000
	CLK = 1'b0;
    #10000; //15220000
	CLK = 1'b1;
    #10000; //15230000
	CLK = 1'b0;
    #10000; //15240000
	CLK = 1'b1;
    #10000; //15250000
	CLK = 1'b0;
    #10000; //15260000
	CLK = 1'b1;
    #10000; //15270000
	CLK = 1'b0;
    #10000; //15280000
	CLK = 1'b1;
    #10000; //15290000
	CLK = 1'b0;
    #10000; //15300000
	CLK = 1'b1;
    #10000; //15310000
	CLK = 1'b0;
    #10000; //15320000
	CLK = 1'b1;
    #10000; //15330000
	CLK = 1'b0;
    #10000; //15340000
	CLK = 1'b1;
    #10000; //15350000
	CLK = 1'b0;
    #10000; //15360000
	CLK = 1'b1;
    #10000; //15370000
	CLK = 1'b0;
    #10000; //15380000
	CLK = 1'b1;
    #10000; //15390000
	CLK = 1'b0;
    #10000; //15400000
	CLK = 1'b1;
    #10000; //15410000
	CLK = 1'b0;
    #10000; //15420000
	CLK = 1'b1;
    #10000; //15430000
	CLK = 1'b0;
    #10000; //15440000
	CLK = 1'b1;
    #10000; //15450000
	CLK = 1'b0;
    #10000; //15460000
	CLK = 1'b1;
    #10000; //15470000
	CLK = 1'b0;
    #10000; //15480000
	CLK = 1'b1;
    #10000; //15490000
	CLK = 1'b0;
    #10000; //15500000
	CLK = 1'b1;
    #10000; //15510000
	CLK = 1'b0;
    #10000; //15520000
	CLK = 1'b1;
    #10000; //15530000
	CLK = 1'b0;
    #10000; //15540000
	CLK = 1'b1;
    #10000; //15550000
	CLK = 1'b0;
    #10000; //15560000
	CLK = 1'b1;
    #10000; //15570000
	CLK = 1'b0;
    #10000; //15580000
	CLK = 1'b1;
    #10000; //15590000
	CLK = 1'b0;
    #10000; //15600000
	CLK = 1'b1;
    #10000; //15610000
	CLK = 1'b0;
    #10000; //15620000
	CLK = 1'b1;
    #10000; //15630000
	CLK = 1'b0;
    #10000; //15640000
	CLK = 1'b1;
    #10000; //15650000
	CLK = 1'b0;
    #10000; //15660000
	CLK = 1'b1;
    #10000; //15670000
	CLK = 1'b0;
    #10000; //15680000
	CLK = 1'b1;
    #10000; //15690000
	CLK = 1'b0;
    #10000; //15700000
	CLK = 1'b1;
    #10000; //15710000
	CLK = 1'b0;
    #10000; //15720000
	CLK = 1'b1;
    #10000; //15730000
	CLK = 1'b0;
    #10000; //15740000
	CLK = 1'b1;
    #10000; //15750000
	CLK = 1'b0;
    #10000; //15760000
	CLK = 1'b1;
    #10000; //15770000
	CLK = 1'b0;
    #10000; //15780000
	CLK = 1'b1;
    #10000; //15790000
	CLK = 1'b0;
    #10000; //15800000
	CLK = 1'b1;
    #10000; //15810000
	CLK = 1'b0;
    #10000; //15820000
	CLK = 1'b1;
    #10000; //15830000
	CLK = 1'b0;
    #10000; //15840000
	CLK = 1'b1;
    #10000; //15850000
	CLK = 1'b0;
    #10000; //15860000
	CLK = 1'b1;
    #10000; //15870000
	CLK = 1'b0;
    #10000; //15880000
	CLK = 1'b1;
    #10000; //15890000
	CLK = 1'b0;
    #10000; //15900000
	CLK = 1'b1;
    #10000; //15910000
	CLK = 1'b0;
    #10000; //15920000
end // end of stimulus process
	



endmodule
