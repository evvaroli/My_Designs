--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:              4:52 PM, 4/19/99 *
--* Tested entity name:                                 Latch *
--* File name contains tested entity: $dsn\src\Devices\Behavior\Latch.vhd *
--*************************************************************

library ieee;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity latch_tb is
end latch_tb;

architecture TB_ARCHITECTURE of latch_tb is
	-- Component declaration of the tested unit
	component Latch
	port(
		INP : in std_logic_vector(7 downto 0);
		OUTP : out std_logic_vector(7 downto 0);
		CLK : in std_logic );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal INP : std_logic_vector(7 downto 0);
	signal CLK : std_logic;
	-- Observed signals - signals mapped to the output ports of tested entity
	signal OUTP : std_logic_vector(7 downto 0);

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : Latch
		port map
			(INP => INP,
			OUTP => OUTP,
			CLK => CLK );

	--Below VHDL code is an inserted .\compile\latch.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

	INP <= "00000000";
	CLK <= '0';
    wait for 400 ns; --0 ps
	INP <= "00000001";
    wait for 100 ns; --400 ns
	CLK <= '1';
    wait for 300 ns; --500 ns
	INP <= "00000010";
	CLK <= '0';
    wait for 400 ns; --800 ns
	INP <= "00000011";
    wait for 100 ns; --1200 ns
	CLK <= '1';
    wait for 300 ns; --1300 ns
	INP <= "00000100";
    wait for 300 ns; --1600 ns
	CLK <= '0';
    wait for 100 ns; --1900 ns
	INP <= "00000101";
    wait for 100 ns; --2 us
	CLK <= '1';
    wait for 100 ns; --2100 ns
	CLK <= '0';
    wait for 200 ns; --2200 ns
	INP <= "00000110";
    wait for 100 ns; --2400 ns
--	end of stimulus events
	wait;
end process; -- end of stimulus process
	



	-- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_Latch of latch_tb is
	for TB_ARCHITECTURE
		for UUT : Latch
			use entity work.Latch(Latch);
		end for;
	end for;
end TESTBENCH_FOR_Latch;

