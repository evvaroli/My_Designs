// (c) Aldec, Inc.
// All rights reserved.
//
// Last modified: $Date: 2009-09-03 16:57:08 +0200 (Thu, 03 Sep 2009) $
// $Revision: 121928 $


// ROM : 256 8-bit words - multiplication with c1=c5=2 coefficient
module rom_rtl_c1c5(
				input [7:0] addr,
				output reg [15:0] data
				);

always @(addr)
begin
	case (addr)
		8'd0   : data = 'd0;
		8'd1   : data = 'd2;
		8'd2   : data = 'd4;
		8'd3   : data = 'd6;
		8'd4   : data = 'd8;
		8'd5   : data = 'd10;
		8'd6   : data = 'd12;
		8'd7   : data = 'd14;
		8'd8   : data = 'd16;
		8'd9   : data = 'd18;
		8'd10  : data = 'd20;
		8'd11  : data = 'd22;
		8'd12  : data = 'd24;
		8'd13  : data = 'd26;
		8'd14  : data = 'd28;
		8'd15  : data = 'd30;
		8'd16  : data = 'd32;
		8'd17  : data = 'd34;
		8'd18  : data = 'd36;
		8'd19  : data = 'd38;
		8'd20  : data = 'd40;
		8'd21  : data = 'd42;
		8'd22  : data = 'd44;
		8'd23  : data = 'd46;
		8'd24  : data = 'd48;
		8'd25  : data = 'd50;
		8'd26  : data = 'd52;
		8'd27  : data = 'd54;
		8'd28  : data = 'd56;
		8'd29  : data = 'd58;
		8'd30  : data = 'd60;
		8'd31  : data = 'd62;
		8'd32  : data = 'd64;
		8'd33  : data = 'd66;
		8'd34  : data = 'd68;
		8'd35  : data = 'd70;
		8'd36  : data = 'd72;
		8'd37  : data = 'd74;
		8'd38  : data = 'd76;
		8'd39  : data = 'd78;
		8'd40  : data = 'd80;
		8'd41  : data = 'd82;
		8'd42  : data = 'd84;
		8'd43  : data = 'd86;
		8'd44  : data = 'd88;
		8'd45  : data = 'd90;
		8'd46  : data = 'd92;
		8'd47  : data = 'd94;
		8'd48  : data = 'd96;
		8'd49  : data = 'd98;
		8'd50  : data = 'd100;
		8'd51  : data = 'd102;
		8'd52  : data = 'd104;
		8'd53  : data = 'd106;
		8'd54  : data = 'd108;
		8'd55  : data = 'd110;
		8'd56  : data = 'd112;
		8'd57  : data = 'd114;
		8'd58  : data = 'd116;
		8'd59  : data = 'd118;
		8'd60  : data = 'd120;
		8'd61  : data = 'd122;
		8'd62  : data = 'd124;
		8'd63  : data = 'd126;
		8'd64  : data = 'd128;
		8'd65  : data = 'd130;
		8'd66  : data = 'd132;
		8'd67  : data = 'd134;
		8'd68  : data = 'd136;
		8'd69  : data = 'd138;
		8'd70  : data = 'd140;
		8'd71  : data = 'd142;
		8'd72  : data = 'd144;
		8'd73  : data = 'd146;
		8'd74  : data = 'd148;
		8'd75  : data = 'd150;
		8'd76  : data = 'd152;
		8'd77  : data = 'd154;
		8'd78  : data = 'd156;
		8'd79  : data = 'd158;
		8'd80  : data = 'd160;
		8'd81  : data = 'd162;
		8'd82  : data = 'd164;
		8'd83  : data = 'd166;
		8'd84  : data = 'd168;
		8'd85  : data = 'd170;
		8'd86  : data = 'd172;
		8'd87  : data = 'd174;
		8'd88  : data = 'd176;
		8'd89  : data = 'd178;
		8'd90  : data = 'd180;
		8'd91  : data = 'd182;
		8'd92  : data = 'd184;
		8'd93  : data = 'd186;
		8'd94  : data = 'd188;
		8'd95  : data = 'd190;
		8'd96  : data = 'd192;
		8'd97  : data = 'd194;
		8'd98  : data = 'd196;
		8'd99  : data = 'd198;
		8'd100 : data = 'd200;
		8'd101 : data = 'd202;
		8'd102 : data = 'd204;
		8'd103 : data = 'd206;
		8'd104 : data = 'd208;
		8'd105 : data = 'd210;
		8'd106 : data = 'd212;
		8'd107 : data = 'd214;
		8'd108 : data = 'd216;
		8'd109 : data = 'd218;
		8'd110 : data = 'd220;
		8'd111 : data = 'd222;
		8'd112 : data = 'd224;
		8'd113 : data = 'd226;
		8'd114 : data = 'd228;
		8'd115 : data = 'd230;
		8'd116 : data = 'd232;
		8'd117 : data = 'd234;
		8'd118 : data = 'd236;
		8'd119 : data = 'd238;
		8'd120 : data = 'd240;
		8'd121 : data = 'd242;
		8'd122 : data = 'd244;
		8'd123 : data = 'd246;
		8'd124 : data = 'd248;
		8'd125 : data = 'd250;
		8'd126 : data = 'd252;
		8'd127 : data = 'd254;
		8'd128 : data = 'd256;
		8'd129 : data = 'd258;
		8'd130 : data = 'd260;
		8'd131 : data = 'd262;
		8'd132 : data = 'd264;
		8'd133 : data = 'd266;
		8'd134 : data = 'd268;
		8'd135 : data = 'd270;
		8'd136 : data = 'd272;
		8'd137 : data = 'd274;
		8'd138 : data = 'd276;
		8'd139 : data = 'd278;
		8'd140 : data = 'd280;
		8'd141 : data = 'd282;
		8'd142 : data = 'd284;
		8'd143 : data = 'd286;
		8'd144 : data = 'd288;
		8'd145 : data = 'd290;
		8'd146 : data = 'd292;
		8'd147 : data = 'd294;
		8'd148 : data = 'd296;
		8'd149 : data = 'd298;
		8'd150 : data = 'd300;
		8'd151 : data = 'd302;
		8'd152 : data = 'd304;
		8'd153 : data = 'd306;
		8'd154 : data = 'd308;
		8'd155 : data = 'd310;
		8'd156 : data = 'd312;
		8'd157 : data = 'd314;
		8'd158 : data = 'd316;
		8'd159 : data = 'd318;
		8'd160 : data = 'd320;
		8'd161 : data = 'd322;
		8'd162 : data = 'd324;
		8'd163 : data = 'd326;
		8'd164 : data = 'd328;
		8'd165 : data = 'd330;
		8'd166 : data = 'd332;
		8'd167 : data = 'd334;
		8'd168 : data = 'd336;
		8'd169 : data = 'd338;
		8'd170 : data = 'd340;
		8'd171 : data = 'd342;
		8'd172 : data = 'd344;
		8'd173 : data = 'd346;
		8'd174 : data = 'd348;
		8'd175 : data = 'd350;
		8'd176 : data = 'd352;
		8'd177 : data = 'd354;
		8'd178 : data = 'd356;
		8'd179 : data = 'd358;
		8'd180 : data = 'd360;
		8'd181 : data = 'd362;
		8'd182 : data = 'd364;
		8'd183 : data = 'd366;
		8'd184 : data = 'd368;
		8'd185 : data = 'd370;
		8'd186 : data = 'd372;
		8'd187 : data = 'd374;
		8'd188 : data = 'd376;
		8'd189 : data = 'd378;
		8'd190 : data = 'd380;
		8'd191 : data = 'd382;
		8'd192 : data = 'd384;
		8'd193 : data = 'd386;
		8'd194 : data = 'd388;
		8'd195 : data = 'd390;
		8'd196 : data = 'd392;
		8'd197 : data = 'd394;
		8'd198 : data = 'd396;
		8'd199 : data = 'd398;
		8'd200 : data = 'd400;
		8'd201 : data = 'd402;
		8'd202 : data = 'd404;
		8'd203 : data = 'd406;
		8'd204 : data = 'd408;
		8'd205 : data = 'd410;
		8'd206 : data = 'd412;
		8'd207 : data = 'd414;
		8'd208 : data = 'd416;
		8'd209 : data = 'd418;
		8'd210 : data = 'd420;
		8'd211 : data = 'd422;
		8'd212 : data = 'd424;
		8'd213 : data = 'd426;
		8'd214 : data = 'd428;
		8'd215 : data = 'd430;
		8'd216 : data = 'd432;
		8'd217 : data = 'd434;
		8'd218 : data = 'd436;
		8'd219 : data = 'd438;
		8'd220 : data = 'd440;
		8'd221 : data = 'd442;
		8'd222 : data = 'd444;
		8'd223 : data = 'd446;
		8'd224 : data = 'd448;
		8'd225 : data = 'd450;
		8'd226 : data = 'd452;
		8'd227 : data = 'd454;
		8'd228 : data = 'd456;
		8'd229 : data = 'd458;
		8'd230 : data = 'd460;
		8'd231 : data = 'd462;
		8'd232 : data = 'd464;
		8'd233 : data = 'd466;
		8'd234 : data = 'd468;
		8'd235 : data = 'd470;
		8'd236 : data = 'd472;
		8'd237 : data = 'd474;
		8'd238 : data = 'd476;
		8'd239 : data = 'd478;
		8'd240 : data = 'd480;
		8'd241 : data = 'd482;
		8'd242 : data = 'd484;
		8'd243 : data = 'd486;
		8'd244 : data = 'd488;
		8'd245 : data = 'd490;
		8'd246 : data = 'd492;
		8'd247 : data = 'd494;
		8'd248 : data = 'd496;
		8'd249 : data = 'd498;
		8'd250 : data = 'd500;
		8'd251 : data = 'd502;
		8'd252 : data = 'd504;
		8'd253 : data = 'd506;
		8'd254 : data = 'd508;
		8'd255 : data = 'd510;
	endcase
end

endmodule
