
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity tank_sprite2 is
	port (
		angle: in STD_LOGIC_VECTOR (1 downto 0);
		addr: in STD_LOGIC_VECTOR (5 downto 0);
		M: out STD_LOGIC_VECTOR (0 to 31)
		);
end tank_sprite2;

architecture tank_sprite2 of tank_sprite2 is
	type rom_array is array (NATURAL range <>)  
	of STD_LOGIC_VECTOR (0 to 31);
	constant rom1: rom_array := (
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000011111110000000000000",
	"00000000001111111111000000000000",
	"00000000011111111111000000000000",
	"00000000011111111111000000000000",
	"00011111011111111111011111110110",
	"01110000011100000000011111110110",
	"01101111010011111111011111110110",
	"00001111001111111111101111110000",
	"00001111011111111111100000000000",
	"00000000011111111111110000000000",
	"00001111011111111111110011110000",
	"00000000000111111111000011110000",
	"00000000000011000000000011110000",
	"00011111100000111110000000000000",
	"01111111101110010000111111110000",
	"01100100001110101110111111111000",
	"01111011110000000000000100001000",
	"01111011111111111111111011110000",
	"01111011111111111111111011111000",
	"01111011111111111111111011111000",
	"00000000000000000000000000000000",
	"01000000000000000000000000000000",
	"00000000000000000000000000010000",
	"00101101101101101101101100100000",
	"00010110110110110110110110000000",
	"00000000000000000000000000000000"
	);
	constant rom2: rom_array := (
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000011111110000000001100",
	"00000000001111111111000000101100",
	"00000000011111111111000011100110",
	"00000000011111111111001111110110",
	"00011111011111111111011111110000",
	"01110000011100000000011111100000",
	"01101111010011111111011110000000",
	"00001111001111111111101001110000",
	"00001111011111111111100000000000",
	"00000000011111111111110000000000",
	"00001111011111111111110011110000",
	"00000000000111111111000011110000",
	"00000000000011000000000011110000",
	"00011111100000111110000000000000",
	"01111111101110010000111111110000",
	"01100100001110101110111111111000",
	"01111011110000000000000100001000",
	"01111011111111111111111011110000",
	"01111011111111111111111011111000",
	"01111011111111111111111011111000",
	"00000000000000000000000000000000",
	"01000000000000000000000000000000",
	"00000000000000000000000000010000",
	"00101101101101101101101100100000",
	"00010110110110110110110110000000",
	"00000000000000000000000000000000"
	);
	constant rom3: rom_array := (
	"00000000000000000000000000000000",
	"00000000000000000000000000010000",
	"00000000000000000000000000111000",
	"00000000000011111110000010011100",
	"00000000001111111111000111001000",
	"00000000011111111111001111100000",
	"00000000011111111111011111110000",
	"00011111011111111111011111100000",
	"01110000011100000000011111000000",
	"01101111010011111111011110000000",
	"00001111001111111111101101110000",
	"00001111011111111111101000000000",
	"00000000011111111111110000000000",
	"00001111011111111111110011110000",
	"00000000000111111111000011110000",
	"00000000000011000000000011110000",
	"00011111100000111110000000000000",
	"01111111101110010000111111110000",
	"01100100001110101110111111111000",
	"01111011110000000000000100001000",
	"01111011111111111111111011110000",
	"01111011111111111111111011111000",
	"01111011111111111111111011111000",
	"00000000000000000000000000000000",
	"01000000000000000000000000000000",
	"00000000000000000000000000010000",
	"00101101101101101101101100100000",
	"00010110110110110110110110000000",
	"00000000000000000000000000000000"
	);
	
begin
	process(addr)
	variable j: integer;				
	begin 
		j := conv_integer(addr);
		if angle = "00" then
			M <= rom1(j);
		elsif angle = "11" then
			M <= rom3(j);
		else
			M <= rom2(j);
		end if;
	end process; 
end tank_sprite2;