// (c) Aldec, Inc.
// All rights reserved.
//
// Last modified: $Date: 2011-08-30 13:31:23 +0200 (Tue, 30 Aug 2011) $
// $Revision: 180634 $


// ROM : 256 8-bit words - multiplication with c2=c4=4 coefficient
module rom_rtl_c2c4(
				input [7:0] addr,
				output reg [15:0] data
				);

always @(addr)
begin
	case (addr)
		8'd0   : data = 'd0;
		8'd1   : data = 'd4;
		8'd2   : data = 'd8;
		8'd3   : data = 'd12;
		8'd4   : data = 'd16;
		8'd5   : data = 'd20;
		8'd6   : data = 'd24;
		8'd7   : data = 'd28;
		8'd8   : data = 'd32;
		8'd9   : data = 'd36;
		8'd10  : data = 'd40;
		8'd11  : data = 'd44;
		8'd12  : data = 'd48;
		8'd13  : data = 'd52;
		8'd14  : data = 'd56;
		8'd15  : data = 'd60;
		8'd16  : data = 'd64;
		8'd17  : data = 'd68;
		8'd18  : data = 'd72;
		8'd19  : data = 'd76;
		8'd20  : data = 'd80;
		8'd21  : data = 'd84;
		8'd22  : data = 'd88;
		8'd23  : data = 'd92;
		8'd24  : data = 'd96;
		8'd25  : data = 'd100;
		8'd26  : data = 'd104;
		8'd27  : data = 'd108;
		8'd28  : data = 'd112;
		8'd29  : data = 'd116;
		8'd30  : data = 'd120;
		8'd31  : data = 'd124;
		8'd32  : data = 'd128;
		8'd33  : data = 'd132;
		8'd34  : data = 'd136;
		8'd35  : data = 'd140;
		8'd36  : data = 'd144;
		8'd37  : data = 'd148;
		8'd38  : data = 'd152;
		8'd39  : data = 'd156;
		8'd40  : data = 'd160;
		8'd41  : data = 'd164;
		8'd42  : data = 'd168;
		8'd43  : data = 'd172;
		8'd44  : data = 'd176;
		8'd45  : data = 'd180;
		8'd46  : data = 'd184;
		8'd47  : data = 'd188;
		8'd48  : data = 'd192;
		8'd49  : data = 'd196;
		8'd50  : data = 'd200;
		8'd51  : data = 'd204;
		8'd52  : data = 'd208;
		8'd53  : data = 'd212;
		8'd54  : data = 'd216;
		8'd55  : data = 'd220;
		8'd56  : data = 'd224;
		8'd57  : data = 'd228;
		8'd58  : data = 'd232;
		8'd59  : data = 'd236;
		8'd60  : data = 'd240;
		8'd61  : data = 'd244;
		8'd62  : data = 'd248;
		8'd63  : data = 'd252;
		8'd64  : data = 'd256;
		8'd65  : data = 'd260;
		8'd66  : data = 'd264;
		8'd67  : data = 'd268;
		8'd68  : data = 'd272;
		8'd69  : data = 'd276;
		8'd70  : data = 'd280;
		8'd71  : data = 'd284;
		8'd72  : data = 'd288;
		8'd73  : data = 'd292;
		8'd74  : data = 'd296;
		8'd75  : data = 'd300;
		8'd76  : data = 'd304;
		8'd77  : data = 'd308;
		8'd78  : data = 'd312;
		8'd79  : data = 'd316;
		8'd80  : data = 'd320;
		8'd81  : data = 'd324;
		8'd82  : data = 'd328;
		8'd83  : data = 'd332;
		8'd84  : data = 'd336;
		8'd85  : data = 'd340;
		8'd86  : data = 'd344;
		8'd87  : data = 'd348;
		8'd88  : data = 'd352;
		8'd89  : data = 'd356;
		8'd90  : data = 'd360;
		8'd91  : data = 'd364;
		8'd92  : data = 'd368;
		8'd93  : data = 'd372;
		8'd94  : data = 'd376;
		8'd95  : data = 'd380;
		8'd96  : data = 'd384;
		8'd97  : data = 'd388;
		8'd98  : data = 'd392;
		8'd99  : data = 'd396;
		8'd100 : data = 'd400;
		8'd101 : data = 'd404;
		8'd102 : data = 'd408;
		8'd103 : data = 'd412;
		8'd104 : data = 'd416;
		8'd105 : data = 'd420;
		8'd106 : data = 'd424;
		8'd107 : data = 'd428;
		8'd108 : data = 'd432;
		8'd109 : data = 'd436;
		8'd110 : data = 'd440;
		8'd111 : data = 'd444;
		8'd112 : data = 'd448;
		8'd113 : data = 'd452;
		8'd114 : data = 'd456;
		8'd115 : data = 'd460;
		8'd116 : data = 'd464;
		8'd117 : data = 'd468;
		8'd118 : data = 'd472;
		8'd119 : data = 'd476;
		8'd120 : data = 'd480;
		8'd121 : data = 'd484;
		8'd122 : data = 'd488;
		8'd123 : data = 'd492;
		8'd124 : data = 'd496;
		8'd125 : data = 'd500;
		8'd126 : data = 'd504;
		8'd127 : data = 'd508;
		8'd128 : data = 'd512;
		8'd129 : data = 'd516;
		8'd130 : data = 'd520;
		8'd131 : data = 'd524;
		8'd132 : data = 'd528;
		8'd133 : data = 'd532;
		8'd134 : data = 'd536;
		8'd135 : data = 'd540;
		8'd136 : data = 'd544;
		8'd137 : data = 'd548;
		8'd138 : data = 'd552;
		8'd139 : data = 'd556;
		8'd140 : data = 'd560;
		8'd141 : data = 'd564;
		8'd142 : data = 'd568;
		8'd143 : data = 'd572;
		8'd144 : data = 'd576;
		8'd145 : data = 'd580;
		8'd146 : data = 'd584;
		8'd147 : data = 'd588;
		8'd148 : data = 'd592;
		8'd149 : data = 'd596;
		8'd150 : data = 'd600;
		8'd151 : data = 'd604;
		8'd152 : data = 'd608;
		8'd153 : data = 'd612;
		8'd154 : data = 'd616;
		8'd155 : data = 'd620;
		8'd156 : data = 'd624;
		8'd157 : data = 'd628;
		8'd158 : data = 'd632;
		8'd159 : data = 'd636;
		8'd160 : data = 'd640;
		8'd161 : data = 'd644;
		8'd162 : data = 'd648;
		8'd163 : data = 'd652;
		8'd164 : data = 'd656;
		8'd165 : data = 'd660;
		8'd166 : data = 'd664;
		8'd167 : data = 'd668;
		8'd168 : data = 'd672;
		8'd169 : data = 'd676;
		8'd170 : data = 'd680;
		8'd171 : data = 'd684;
		8'd172 : data = 'd688;
		8'd173 : data = 'd692;
		8'd174 : data = 'd696;
		8'd175 : data = 'd700;
		8'd176 : data = 'd704;
		8'd177 : data = 'd708;
		8'd178 : data = 'd712;
		8'd179 : data = 'd716;
		8'd180 : data = 'd720;
		8'd181 : data = 'd724;
		8'd182 : data = 'd728;
		8'd183 : data = 'd732;
		8'd184 : data = 'd736;
		8'd185 : data = 'd740;
		8'd186 : data = 'd744;
		8'd187 : data = 'd748;
		8'd188 : data = 'd752;
		8'd189 : data = 'd756;
		8'd190 : data = 'd760;
		8'd191 : data = 'd764;
		8'd192 : data = 'd768;
		8'd193 : data = 'd772;
		8'd194 : data = 'd776;
		8'd195 : data = 'd780;
		8'd196 : data = 'd784;
		8'd197 : data = 'd788;
		8'd198 : data = 'd792;
		8'd199 : data = 'd796;
		8'd200 : data = 'd800;
		8'd201 : data = 'd804;
		8'd202 : data = 'd808;
		8'd203 : data = 'd812;
		8'd204 : data = 'd816;
		8'd205 : data = 'd820;
		8'd206 : data = 'd824;
		8'd207 : data = 'd828;
		8'd208 : data = 'd832;
		8'd209 : data = 'd836;
		8'd210 : data = 'd840;
		8'd211 : data = 'd844;
		8'd212 : data = 'd848;
		8'd213 : data = 'd852;
		8'd214 : data = 'd856;
		8'd215 : data = 'd860;
		8'd216 : data = 'd864;
		8'd217 : data = 'd868;
		8'd218 : data = 'd872;
		8'd219 : data = 'd876;
		8'd220 : data = 'd880;
		8'd221 : data = 'd884;
		8'd222 : data = 'd888;
		8'd223 : data = 'd892;
		8'd224 : data = 'd896;
		8'd225 : data = 'd900;
		8'd226 : data = 'd904;
		8'd227 : data = 'd908;
		8'd228 : data = 'd912;
		8'd229 : data = 'd916;
		8'd230 : data = 'd920;
		8'd231 : data = 'd924;
		8'd232 : data = 'd928;
		8'd233 : data = 'd932;
		8'd234 : data = 'd936;
		8'd235 : data = 'd940;
		8'd236 : data = 'd944;
		8'd237 : data = 'd948;
		8'd238 : data = 'd952;
		8'd239 : data = 'd956;
		8'd240 : data = 'd960;
		8'd241 : data = 'd964;
		8'd242 : data = 'd968;
		8'd243 : data = 'd972;
		8'd244 : data = 'd976;
		8'd245 : data = 'd980;
		8'd246 : data = 'd984;
		8'd247 : data = 'd988;
		8'd248 : data = 'd992;
		8'd249 : data = 'd996;
		8'd250 : data = 'd1000;
		8'd251 : data = 'd1004;
		8'd252 : data = 'd1008;
		8'd253 : data = 'd1012;
		8'd254 : data = 'd1016;
		8'd255 : data = 'd1020;
    endcase
end

endmodule
