--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* The configuration file can be used for simulation of      *
--* backannotated structural VHDL files.                      *
--*                                                           *
--* This file was generated on:              8:02 PM, 4/20/99 *
--* Tested entity name:                             A8051_exp *
--* File name contains tested entity: $dsn\compile\A8051_exp.vhd *
--*************************************************************

configuration POST_SYNTH_FOR_A8051_exp of a8051_exp_tb is
	for TB_ARCHITECTURE
		for UUT : A8051_exp
			use entity work.A8051_exp (A8051_exp);
				for A8051_exp
					for U1: FPGA
						use entity work.FPGA (beh);
					end for	;
				end for;
		end for;
	end for;
end POST_SYNTH_FOR_A8051_exp;

