
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity player12 is
	port (
		winner: in STD_LOGIC_VECTOR(1 downto 0);
		addr: in STD_LOGIC_VECTOR (6 downto 0); --8bit if WINS added
		M: out STD_LOGIC_VECTOR (0 to 41)
		);
end player12;

architecture player12 of player12 is
	type rom_array is array (NATURAL range <>)
	of STD_LOGIC_VECTOR (0 to 41);
	
	type rom_array2 is array (NATURAL range <>)
	of STD_LOGIC_VECTOR (0 to 22); 
	
	--PLAYER1	42
	constant rom1: rom_array:= (
		"111100100000011100100010111110111100001100",
		"100010100000100010100010100000100010010100",
		"100010100000100010100010100000100010000100",
		"111100100000111110010100111110111100000100",
		"100000100000100010001000100000101000000100",
		"100000100000100010001000100000100100000100",
		"100000111110100010001000111110100010011111"
	);	  
	--PLAYER2
	constant rom2: rom_array := (
		"111100100000011100100010111110111100001110",
		"100010100000100010100010100000100010010001",
		"100010100000100010100010100000100010000001",
		"111100100000111110010100111111111100000110",
		"100000100000100010001000100000101000001000",
		"100000100000100010001000100000100100010000",
		"100000111110100010001000111111100010011111"
	);	 
	--WINS		23
	constant rom3: rom_array2 := (
		"10101011111010001001111",
		"10101000100011001010000",
		"10101000100010101010000",
		"10101000100010011001110",
		"10101000100010001000001",
		"10101000100010001000001",
		"01010011111010001011110"
	);
begin
	process(addr)
		variable j: integer;	
	begin
		j := conv_integer(addr);
			M <= rom1(j);
	end process; 
end player12;