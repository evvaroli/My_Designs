
module top;

	reg p;

	inst #("abc") ii0(p);

endmodule
