package maths_class is

  subtype single is real range -1.0E38 to 1.0E38;
  subtype double is real;

end maths_class;
